XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v�LB�O�?�DU;�{��gq�$ࢩ9�S�ǆ�i��:�?��6Մ��͢68?��'����;}Y#�MA�]���C|���"͜�cn�I�
�P9ZZe��\�v�p���RBE翞w"�D�S�A	�Ƞڪ/@����i���Ҧ.�z�R�Ԅ��Ý�+{C�Gp۟���Q�C�U��<G�$H���:���E4Ú|h�7�^xD$�T}K4�^�嘭��sh���Z!�W�U�P�WS\�Ud���,����I�G����^���mI��L\E�+�W0���\I����"(ƾ�!�~�G<��hX[kk��E毛�8�Ȫ[�Y���$���Yb����W�pL��@���b�u��BM\r�wӲ�R6u�N�G'�zC�_hr�Ll�r���XoL@���*V�0h�F�>�B�wN��@Qz�t�P�ȡ�'JY%]���x����-�6�z��?��5N��	Ǳ����e;��p��ri��Vl͇0�r�z�u{�IR:���R8�N_����ad��(8#��~���i��Y�|��wu���L{��']�8����f�S����	h5��x��w�kpb�	��e)Z@�ĺ��8[�*iɂRn���g��'.SQ7ZBE��-���T����1���x�y�.��}��]𦩡���"b)�)����Nq2/��Ǖ7����5�1��2��'���R�	�����2��<�6K�>�3	ۗ�z!m��sy�5�w�1���4W�NXlxVHYEB    39de    1170��CuO��,o�t<}��qKV�U���Ox���ų���ku��u�ڪ$�jr��]M� ty����Jߓ�-�b�������Ż(/|��RU6ׁ���!(ݐf��W6��Dx���s�VU�o�_t�����~DiS-��=t�eZ����"Ŭ2���ҩr�@r?�˳�FR���z��(n`U�2w��L��������J�<Ta��&��<;��/"�QE֜��U.������v�/��,IQ1����S�n�<dO����L^c�V4�B�4�-�W�J>,c&Zg+�M%yz�&ЩN�d����<֫s,�Y'��t�����R.�or@���<6�  ~P#Wժ��ʛ� �A�N;ŜI�庾��>m�}�(Tk���j���'DO��=��ƀƯ���߇cx�h1��am&�R4���;�^�Q���8�!ˌdp��c)A�e�Z2��/9�}���f�=3>�#����g
c�n�$o�c[D��qEۍ�j��0���������y2V�w�$c�?ɰ|d��[G��B�J��,�:��b��
��.�i-�� ǵ*<|@��#���TGˡ��}���n�������W�_y�� �*<�_׸; ����%ZLi��WY�ik�@�*�<1�
����M�_ l�2ho��};pyU���gO;@�HU{�3�M
c�.��� T|s92���1ze��������C���~{��h�,�ջ�풩�s���&k��YUc�G$�*�[O9�BD�s�mEb��6r��!�/}���u��Jz��~�DB!�2��p�L�SL�?MJ����t0��.m��.�#=N���}'c1-� $G�♿f���O���U��K6X�"Tƶ}Φ�p�e���bN #X�X� }�ni���.B݃ |<e�����9�1��а1Ĭ��c'V�2i��0n;C���7����ᢆGN�$&��e�b������p_����Eb�`dJ�I�0h���b��%nf	Ih�]�.?�p'�~�Ouo7��1' `�-�+�ݗ�O��"�t��	����T� �}|mB)�;2��_A�P��ʁ�|�����8�Mۨ��3;�~g�,���_���_��7�U�lw���k��(ݜ��e<�	GSj6&(�>{%;{w��R	�/��dT�~�p[L�'�@����Z�<[3�YuE��}K�����OC����`އuF���Ч?8 �l𗵺zlC�r�ͥo��q`kuf�2Z�����L
���9\�*��dx+@W�`V�+�U5l�y�صܚ��C�o��=�m2!��;�4T��E�w)cX*#� �&ꞙ�������yt,�����+�nZ4�B�l���׳�zWK��**nB�Q��>zX�s����is����h2J����i��A��6��m2������4�:���b��H�wSۿ�a��zռ�+e���E�Alp�E��w�	@(�9�g��Y�Ap�@��X����[I(v�Kv';��o�]����.�o��:�l�ZjVc�.7=V�'x��$�;�M�P���SO�BĔzuh�\���|����6��<����t�ah�Jx�,۩'�{`�R�xm1�
�柙9Jb(��/��.x�(���x��OgƬAe��[ѫʹ!��5E߭~��w4��>�Isݾn�E��2ze7��=)��m�We���+{TW-�4oy��{bU�oH:�Ou2:Z^}?��pG"�dՁM���a f���8^�-�S�櫦�����3Ќ����O�U2&�w ���r*��o����,��!R��8���1���K�g�������S�=c�Q��=���0r~?��i�Ѧv8�SW~O��;i���l��y�&��Qh��F��23vJIFiK$*�g)��=i���(��;C��` ��Dx�Tq��J_Z�\;�S�L���<ñ�^a�u��ٸ�\|2�l��J�����A�o*
H�,x����R����E��K+��/�N�C��4�a"ǯK /|����mqa�46X��o�c�d.�j?)�Ţ�+��ƭ�nd&�H�uֻ�b��p��2D�D�e�ʱ!t�O����uqses�|0�g ����{D$�6�<����i��d��SD�0X�x���"$^K���n��m��}�#�Ж� tڎ����^A�X�������������X�� C�R{ƞ#��s��"#����Z��]T��x���B�8�'��[,y�׃f�����@�L��M�!Ъ5�<�`���eO�z��n�k�����G����L�D�<ۄ�{K��o����JV #��5�9�Ox�YV>	ok�Ќ��_F�6�i����c�b�x�&v|�]X$�焟l�c���hD�
�كK¼}�%�u�`�znv�#���ґ`� ��?�j;����yXX>���s�=��5m�O")?ˁ+J*n�Mۼ��j8oo������ti���lS�������b�7�C����?j���T���⟩K�A�{����1�{���0�/X��T�7�L�)d�b����g�i��p�T��B� Nb!��Q�G6�]�7f�%��ح4��zt�-,��ݟJ(d����a����iK�x���1��;���iRr!r�TKG��sh�k-�|]�Y�t�RP1-�1�E��,)��IK5~��~P"�795^�18>��	Ĵg�yQ����;�b�&lRX��Y�u��el��A�a�7�}��&K���� 24�Ӏp�����~rL��\Rt�
n���s�;�Rn� ��z��3���B�Β)B+&0��B�_nWdꐨ���>�Wo��Й�䟀�fcC�S�bw��{!>�5�3���.CV�;��W��*�r��D�^�(C��9c"��<�}?u�"�K���zo�}��d1���&�P�jb����^\ʴ~|M;b��A�d�r���DG�e,�w�a׺2�����FMIW�4����?v
�:h��s�
p�rm�q�c|�,�6+O�g{_�H�OG�~����J\�z�a`І�$V�f�L��N�t�W�D�C�ca|��$���
k�?�I�Ds#5ъ� #,v�VK�%@�J%󝲚n��V(������\R=.i�P��`U����r�7cBQ�z�/j�;��t|�?��\����5P8�罹\Y�'�K��`ÝO2y��;�o�]�l-�']�Ӊ�k��ik��?g��6[�2���S49�K	�g� k�t�	g�T)��ApA�j����ĭ դ�4�N���f�j����E���S��Gڛ+�/1k�؝hP���7Z4��J����/>2 n'#9��C�O����H��߸�7
&g8��������ѩ�`Lt���9��qPZ�#�UqX�;�r ;�jV�-nձ��0Ԓq[��{A&�~��y@ik/�/��9gD���%�{4���C�v�L�TLQ�	`���������i�*Z+gJ��A��J��k�X��I⑫�*C�-��$]�P�[�n� �
i��T��r�/B�>�<��׵䡡�(n��y���#!v&��_ř�B��	�� QT{�w��L	�49��Iv�ګ���n崴4&�h�s	 $f�I:� ��p����x3��J����Ĺ��L�rq�i��9B�rL�Z�F�l� @wS��ϻ��!e�H��V[��@=��D�C������n�cua�K%�!�R`+<�?F��tJk(�9Ĥ�,��0�I�e<$	Pˏ'ꄧ�it�Y���u�E漛��`,J~3_�K���4�SJ,dW*[���G���{k��Y��#!�iL�^��������W�Q���a,�u��ӧ�iF��yS���Xa��rWj�rױ�  ��n�!(����0"�?}74E�v��6�p�Z@f�0������-œU�U�� 1�^��E��cj��5�a&����?@��_�:��P����>�x`���i�I@&�Ra�8��WA��Cg���*p7{Y'1 ��D�p=�|x��v���p�pwM,y� �!�Ca����������-*W��ԓ6-k�$�Z�0��
M-�C��v�lYѳ��x^��Qp�8B�l-��0�{�|u�)�ۙۧ�*,��Cn���K,�7X��gB-�s6%f�.a<�ǖڙl�Z���������)��%(��H	K~t�`5�V�O	8�PD��?�Te �C!�����������@Z�q�����z��狃$%�)���&W�\���כ#��n��M��P�Է`���.r��'Eb���C%��Y��Zr��9�V�s5	��� ��^P3ϔ�fE���FX��Y���U�}�����7��m蓙|�x