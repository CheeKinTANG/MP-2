XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����*=��s�]��\.y��*�ћ������`2�Կ,�8הn�r��p�N_Ų>��RqH��� y�.0�z*Y�{(�<.�V	v9������/|������L7k������`K��A��s�ݏ��֧����~^.����AT�إZ5?]T˳8$����ٶ�P�W��� �[D��}]�d (�����E��o��S����v��O�Jq���	
�мC
`"3�|b�$�5�j@,x�7&��!�l�	�y��=�D�
�!��[��q�e���W�%��Z�o���{Xk1����$7��ا� ���	<���|V9&$T�9��{����;� ��&���1Q�*Aa�{l=p���{�M�a~�&���5��_��T�h�I9��	���I�W;#9-#�$�R?A�i�c��B���Ҷ�����xo��NS�?s�K��߈�`�P_�N'���U��:�a�Ic�8�d���oڜ����	��A�����܏��ƿk��l(A���24!`���%�V@_#%2П���!����F(��ؓMB�t���K�d�;Z�<��Wq{@0�w���y褵�؀�$:�a;P\����3����N�%Y�5��@�|ʻ`8#�Q@5����k,�}-Pr$~��o=g.E&�H�S%q����%?��W��[��O��!��}���z�YV-���WQ5ޜ�eIh�T�w|�@"o4���gع��߶�T�S�[Hm��yXlxVHYEB    3fdc    1160[�"�Z�e�D�}&���,2ȹ�M�0#��Ɂe ����3���p���g�1�[;�o�p�چ����Ar�������5Wh^qN����.�h1�Z��^(aB~;�k-g�_�Z�h��'�Y�w֏���Q�|�O['	��7 q�կb=P�J���>p$7��?%�p3�� g��;�j��+�Y�e����|�ʜ��`���Y���G˄��E�,Qt�ʠ�cmC�8!Z�<KsНj

��<K�vD��]����k	�)�Δ:+��h��g��J��[�d1��&��Uࢗ�D��Cj�x�^d�1��Х�n
tCy8ypA���|0�I��P��cp/�6W��-pFg��֞Vr�y�� �z�ߝf�*j�
�+b��]���
aV�d�eP����vb+ܧ�j8���Hd��x7IX��g���k; :�*z�d����)�"83V�t l �o���1��s�"��R�9,�n0���s���S ��Z�R��3��m��(g�����h�J4�F+��.8-�/�CQn�N�dc�ͨ�
����gE9��=���IV�O��?�k�R�K��	���k���J!_��58�KNZ$N^Y�U8����FR%Iyq�V�!7�ZNHv��&���)dBJ��Tô�(>���T�J�B#:��BOZܻ�.Q/����э�EG��BSw��BR_M:V`�ӸA�P�$��F=Hx����뉤VY�*h�����DVU�|���ʖ&���� >�#�e��	H�[O�@k�T�A��d\8l
���:F�FK�J�H]M8?�|)��0�K��#㎁�`-���`y`�sB�%$��g��������<��c]��͗s6s�*��ׄsO�@���B&,Gf���V��x���X��� _V���q�3���1�G0¬w^]xm}۵�=EOr?�	&>�*�F�Q����7��4禊<��j~��p�Ƨ��|�?�.����/��DYqC�}�:���t�ۑymF�a��r!m���ׇ5�B�$~Y��|$n�t�+�en����ۡH�k��Bd�l���/[���w+ f���uwð &^��^4���݅��8w�/+)�z.��5,4�bڒP�w�>/���k<�r��-�����B�g����Ȩ,�Q��	�x�����ߗ����m/ɨ�`�>��7���O�����jBA�&o�fg�����`�紨��CdW�D%0*��4�Ig藚��LvYwl}��ݹB(��[0�o9�HC��#𬍸��`���XB�w����f�Ig�"�@4�5���n�enָ8Vx*�Gp�����~����:V\O���y�*���>��y�>G���d1�
�����H�Z�_Dt *�%�$�'-�n���T�9�K8X�ΊO++��|�XOZ��9���|�E"��۲�zlB4�4	��Ẕ�V���5&֩�gQ��G �G�o�h���!�������h�(�6��ozV#��a�����׏.��>RݲS[4�_�h�މ��Z�^�1�9cP�T?���%�v��ѻ���T�'I�m�s�S�����uv�wQ�]�����[n�敫�E�rTNص���ѝ���zڽ0�)2oda��/��1#]7�h%Q���#���Q"��ë�㫅#�.�]E7&�y�����R�²:m`���)�����sp��e�j��N*�p��vE(�|��G$�H ���I�(���{������5+#�[!H΁3>\�t�V���=x1|cۤ ��˳N�{(C��2!g���y���������?i�{Cϫ��?�=Z�ג�񠤴P�r�e|=c]R��q��H��sjo�oq۴+�VOӘÚ�� ѵۧAB�%�
@̋�1Ix�1\/!Gh��SI0�3L腭Y(@I�Z�\ 6�fݞ��UG�h@��. ?J�f�h�¾(���`�ޛC�Ij�"]+���Ul�(�3�{�@*]��y��W�e�ig��b�|��!g�4�������3>�q�Θ��._�����k��?~�E�Zp�	��汌h�G��`3�J8ڟ��A 7Y��?�g��tcXu�_�!,�e?S���~�)YM���,7�߿F��	��A7xdq�T
k��s#l��R�Ь�Y�9����E������}�ܔ��c��A^�0$�/��û��?D��A2�r?�[���6�߱k|;.g.�J���A�3��1��XfV�Q�!�B�/z�6�*G��N�A�B��.j�lwR�?7R�n�:l�8����#�A6�K����$X��W��FkOf�l����8~����nB��.o<��8@�����S�-nM��O���gf�'&��;��Z�'��9�L�M���Pߊ:�����J�^{�2Η�o��u�~���K����f;V��ʗMTn�m� ����;+c �ܡ{V�J��Kʒ�|�$�#q.2yYHA-S���f�M5�"��^�c{�N�U:࢘����ƒ$����eЬ5y�3��,�g�R)���<�%�V�����~}l�,��N|~���|Oj�x��������%����?�c����H(7\����l��-�%�7�CI}�Y^�di̆���R\�h�-[5>��3il�jg�,*�D��W��{Gt��$�G;��]B����9�#fhı2�X#�;�k�t��*�vw�z��B6�J/$���wzv�A	�;e�fȔ�&�1+��K��.�b9����W� a:���ǲ�YsD=��{��-�jn\-���.�Qo��^}d~�,��Vu�#�p��z�
H�pF�� ���7^�o�r����E����� hS��UBo)m�Q/l�U^��{�kyP��M�=�C��ۂ��]74�����fd�w�vp���9�=�j�`J��~ D��%���d�W�+�^��!�y�#*���"��_)|P�ND���}�2����{��G~���D��rGL9�oYn�
#���w:�i G���S�aE��BU.��^(O�q�����&���%���>��m�l�)x'3�(M�ⓁO��ʙ�[��������I%�f�E���X���J�)�C����Qj휰��]��;��&�z��Wd۵�p_�~i]�5�joq��L�I@U0�i�3S$D��O�S��$md����m�ȃg3Y跤)5��@����K�$|"��c	���;���Z)UoU�翄mՖ�p%ڌ��y�EF5�r��9"2yM9�?�pN���'4<�]���>��d=��~Df��2�ۚj?O�����������Ҧ���vU���	�.oԋ�!��D$F����֚1ګ쟴P@M�
*�
��},w�/FE����b<�G���[o�S="y�)u���-�"��x�C#q�=�*�t>�=�ó�Y.��#A�ы��zE��%!�
�;וt�h1�n�t���Q�B�Ea�Z��z�*c����pv�6���ku7�T��b���l�ue������c���䃐��xtBǮ�P�v�K�<|�;��:A�gI�W�N,�}� .qZ�ӟahk��԰_��د�����q�/z7��/�ⵢ�.Q	"I��v\h;I���"'Q��OI���}<��{�k�����T*����_�)FV��5��(#��s�5��C�����!N��o��F������@��$��	���}���ޢ<Wo3Φ�l�M=~U�m��LQ������)tq��n�IZݮ�a׽j�0��D{7񍨾#���P&=&�L�є�P��8� �;n��v��x����G���9�Y�R�8���uJ{(�^��S�M�d�k_�V�_�Ď:���R�t�̒z	�8�8�f�6Ư��U��Ɋƙ�l�:�{�Y���/����(�19����PH�)u��%g�����H(4hcF�,z
��7D��4���_kt%��댢���H��!�Z�Q�F��7���V
�	/^Ј�'�N�!�K�u�[�t^����	�z�NS����j}\��2�q`�&�Ŋ���W̀/R�T��Xb�ȿVVdܐ�r-,�y὾e�{m�;�@L�}�A#��AG�~;���AkrA:tnx�aJ�f'r�\�~�=�!:ɾ�+{���*��>��m5����Y���2��pȰ�W�5�p$�E��pҿ�Ra�+��j�~�D>�\*��q����tnINqE�n=���2=��j�ڱ6�G욓	X�\(�<f�?��B��}k�
�ե�7Zzűz�����Ԡs*n�#.��$��5h����� ًt 	�p�ǭ���*��Cc��@�\�Z��|G���@�/	|���M^��