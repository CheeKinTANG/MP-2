XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����K����<nȍh����$~���# ��/��?�wцs-����޷�ht�qp��Es��Ȱ���T��x%��)3�!�<)C���)�����ΉNc%�,�!��1�x��ٚB+�\+|D���������t>�R�U!gP�4���į���N{�>�s��͌��%%z$�/���Ev���N�L	�.����g�;C�L�a�K�?�zd/��ؿy��J��k������&շ� q�2��°E��~�;��qEU��f}Kwp���pd�^}h(���Y5�e�n�N#+PL�~�U�t_�%�o�bÏ4p�}����u={�Tي��De�ۄ���t�k�j���.�|3>ˡ$^�%�E{�J�T1G�^��ʺ%I���
mEsˮ�6������H�)L���zd�wL�tI���k�|��R���X�#b�k��j��_Ǣ?�� ����<���L"6_���o�6'�5G��1N<��utc^�`aً`\�%V��b���G��r���ck9�آ�"�\;����k����v�p�p
��t����ޔn^���N'b��EҎ��4���]���Ok�@��=�����o����?��Ɇ���`]��&�]�OC��?1}9�1�	�d�M�I^��3�Y�KoK���E,M2CG|s�M���a1)�;LM��;x{���ޚY��;�|3y6$����`-qoЉ��E��!v�ؼ��R���U���|"ff�v�ut[x0�"��\��Upm�Z�,�!XlxVHYEB    b087    25404����d u�i�g��E�	��7{���ɨ�H��L�&�^��X0��=�p�S����w[�tW���"g��N��{��­�bA���D0��>4�H����3����-V/O�"�{��Ӵ���xvu̒)�,֨�nfjLN�Շ� �ZVo�9�ʁ�;7Ă���b]�6�@��/��sT�3�WQ%��v$�c�Ysc?�G�?�p���1�ŷ�
D���_nV��R�)�t�	�"�F�PR���`Og�C��)���>�XC3�9C�SDL�JO�g��;�U�w ̈́�h�~9=��Y�CdT&8eK7��B��m�z�Η��o$u��}���ĿMR'mҤ��aw|�9�Cv���U{�B����}mJ��G5�md�d7��}p��s��ޮqYs�kj��w<U���O�ᾪOU&�&Ԡ��*�w:�Y~I�Z�Λ���PyA�q�X�whkq�)��&��o�.y�b�!��0.���d������+�/-���n��M��e�{[�O�ͱLI��j����ǁA!.,O��C.u���-�J�c��c��20�3n�bab+�,�)���0%L�^��!�I(�h�sR��^2㆟� �xx;��M��?�mB&��"I�)Z>l��#5���3_F��+>����/������u�:��P���)��
1�n���"Z�� ��#���H&�W�`�WV����U,��r\8Ov>��	���`�r�m�䱁��
_�;�w�b@��Lq�8x��g����|�}\тa�`mE҉��n�`9Mw�yM�O���+�/��tt)jQgDk�
��!�y7���}�X�^���JA���B���$�ѷÛ�p�������I$=vÛ�t,���}�/V@��^�l�HQ����%c3�tr��Ѝ��:;/�[@ ^1��͒6����X��E�1_�h0����蚨���� 51�0�g闀~M4�Pcp64�o&�\�E6V)�=zHai�"/8#��ͱO��?��c�C�G2%kM��I�Hԁ��ۼ��;`U�	ox�Ȍ�
�ŚW��;���H��ä��1�����q���T1dZ���g�O��Wg!}|M��������L��d��a����w�2p�m�-�6��'�\���[}��"���@�HWa7Lw��O8��p�k���&\(/=1\��p[�A��$��ZS{�ay��ئ?���$�[�(gN^�Fʇa�R9��I��<ĳ�V��WŚ5n$G�*D�+i&�9e.��Ь1�p�Ş�\?#�x�>|4}W&e�ic�5���(\�?|�55�	l3�zQaDy�;r5_�Zu��|��	jO!�N5�$+��.�I�Z���k��"��f�+�X���p��n*a�[���p,���7�Ȩ^�I?Β5�3�~ܕ8�k�R�4�ku���x�$�����{�ۘ��z?t��[�������&C&L�K��4�1E+
�(�8���iG�:��sE[��˻|Ɂ5N�Q�j�W����<�L�وO+./g`h������S)�x�$����M�+݃|Mݮ�pƇ��ڰ�ܳygF���6ݍ�6_�c�"��$'R4.8�!�5�\[o7'��j�@��sX�����%}��C���Q��1I�F�^?�:��I�:��`�GĦ�f3�T�C�ћR���|e	F\�D<�=�������q�fB���ǣcf�ӟ�F���E�4�N�!T����P�x�bU�xX�6�J:����`[h�76l��`I0�"T�b	NU��b�+0�x��5M�/Ұ��6Ĝ�W�킟�7�L�HګT�]�S�B��p�/FO���C^#٭�A����TT����*Y�������T�p�{�<�#���/r�pC@#GÏ6���}�}|o���ь#�����g�؆]}����� $�Z�;���U�=���8�B�/k*:�^)��=99�$�߷2:7�"�bZ��2�4!��� ˈK��gg����3V]!�?�m�s�5�>3!�*���*E���c��xիG��ZZs�@݄Y���^4��яg���-�����[��cF�o���Ґt� ��¯�`%5���h��<�~���ø�Z�B��_!Y	6#����P��)4.�����uF�>�����i�n�^��/�	=��������������Uu��x|�6%���dG!�K������ܐ�H��:}Z^�P��h�������7xE�A� !��9�^v����}��IU����$���au����w̬7rS2���U�Rd����kI�\"��{@p���El�Y�)�qgB�u/��-��y笣���G��`{\&-�z�x����\'Jir7|��a�ꛂ��@F������u��"$��ۼ���%l�����k�Qu�u�_c@��K��2Zt,�+����q���a�hH�og�1p�D�����z4�7���aU��gMua�l��Cd���҅$b���q�dnps����'�yFz��x$��9���I�#@�9+_Wď���,�a����$�w-7ti�d�\�9�/���>g+W��J����������C���-;�0��j�� `��$PY��e� ��%˨�%�
T]��W�ao�����v��l�#��}�B')��O�/�ѩ�upO~%�|�u0���䛁�O�V�{"�G����jj�@�\A���2��$��7g���Tb޿)��l3u���N�BW"M��jH��c"-�1W�\��V_xW���Vbʷ2p��"qT����[ۼ��'8�@�ݼ�8h[���*����Gϳj�rKd:�����A�*;�l��A�1ݗ��)]틞k�tEn�r	x�XE"���� �[k.�B��Uy��D�|�
���CHy���DSe<��V:EL�*-���}��[��l��r��2)�x�v��������<��*]�;�Ը.V��HU�fvO����ؘ�n�0v�K�	���N���x���F@����q$���sf`ǵ�Y'�Ff5��HV���]����s�ܬ�m���(�#b��}�yW�0��+�m�i�V�d$;���J�I6%�	kP���X��L�x���>�	Eb}8Z�;�B4J$�z>�R����p� ��=E3�k�}Qw��fn��,��=O�㊃���B~��Z3���K���%u�{TTQ԰�����#���]clD���}�	o��Y�f��ܩ�֣2�n&���2A�?��Z���W����@h� ���C	r,����c��ԧVsȤ��1���%g��R�
��Zq�����9��K,s{%w_��ց2&S\���7Vͨ��l̜��]�O�f�?S�P͹�9\�b��*��&m�ѻۿ�/�ў1�uqFݓ�c���#:C�|N��C@935O����磀��E�6�"pB\�RAn�w��5m�P�*�*6P��3�E{"���f�^3�x��~�R!��A5���,F(S�qt�/FnT�@��DՁ���`G}j�'&I��ᅱ���~?�m|�kQ=��
6��QF��J������5]�2���s��(�@s�?c�BТ]��4�YB�"�[U�$��(,6�Z���=�y�<[�}��dF�ʥ\`��g'|�j�ݶ�ۄ���t�;j����)�l�풎�
,:>R��1/?���C�ݼ8����=q�/�����?��d���zR!�]�?�?\�5�������ǽ �9��,^1};��[� ���G�Q�M c֜~sI�^����-���ckR+���Z���ЄȾ�$�8ߐ�z�A�~�X��C��ܯ����q_���ћ�c؉����5�w^S��TJ��T�����;��&�ߖL������������g�~N���ii�	/� )�? ���4��w?q�ur����A�e���e��ƠdI���7�Z����9x�6�%yGB��Ի��v�b�Ҕ��<��;ǗR��^S���vZ7���>�iZv�]q��;�	MA	��Lt������zo��9.��Yv_�����Ljh�R��n-l�Z���g7��Ȅ�48̎���b����֡.������.�+�V�� ��3@-V��Ϲ�X	�1��(V��һ�b#VJoW��8ҋ�<P,©d�� I�hM�G�X�o�a)��P���l�VPv"P�LA�r¨�� <�iu+�/�M����=�[�!���%\����A���l����V`py�|��L����6"��!�泥�%�	�7BE�D��])H�'y�N��,Ŭ����+�ʋ�:��<eh�X���:�%x�t�4��bq7u=���`	�;^�/L(��l� �E�+Y�k]��|���3)!7��1��O޵��,�mb�����X�L��;��P�r�O=��W��;��.��o#�x��i���b_w��� lZ� ��Ƀ�~�'x����״cz�d���}N��[�0���qY�D�M��L��"�4N����@0^e�&����p�[����5����F_�m#&�ЋS����������b~��+�]n�3�
l#�y�]T殡^ +2$����<����mW$,Ʌ�5�n"�;�ѣ�;�$q�-჊�T.	Wh�U�(.��	���OX��z�Hْ�:ǶO���T�m4�@��m����R��ky��s6YD"�iP�W�Z[ت�y�t��B2A�}<��S��T���y��q'TĊimS�Y����<���(Xt��t�s�l����3��á��EԘ~�u������a�љ��9K�f��gu�"LS���Lkj��-��T�/HH�A�݅i�»�/�6��� ŋ�04C�-5���������鏐h6��2���<q���>��3�	�Ȁ�W��:����n�!��:E���ũX�1�9g�mu3��q@lx��*�EXc��ku�
�a)����<1�#bw$�]z
V��3��1\bk5��uI���6��	��܍c�Qjkv��URuM�F���°��~�i�3��oIϿ��Uk�C���6����%���-j��`Y�)��L����B�ge�7x�t��{�U+I�ؿ�߿e�A@�g{f����N��sE���W��A��E����ek[}|�n����e�6��P���U��c����Mre*"�E� ~t.�G[w���T�������vD�8��}��)=Y��)lY�>qB�I��}1��fm��Q���u���� jؔ���1��w+�˝&m�� �Z-�C� �`�
�"�avyiJ���n�r�Ɛc"K� �N�3�?� ��Y��� 6N��Y`�w�c���f�yg�^њ j�L~T�i����F�賰BP|�*?��	1�p4�(;�o�I�
���	���P�QN��?m<|���L���p`F����w���.��J�F�7\Lg��e���r4H^�~@F:smv��
��XT��k`�L�5��7�O��=-tK�Q� ��b�������(���a�c�-U쓊N���f�Wy��X1>.�����`h�HW�F�L�;%ٞ3�$�>��d���5'S�x^j|�6�"�'�Fb#<1��m�b^N	�Ш������AD����]4�h��L=1����_H ����	��w�w����6�j(wF}k��8��awʛ�&N��c�vv� ݘ
׵~�Lw5#���Ѿ�ҍ�S�A�� �梓��>9b�H�O��<z��9uě����-�h��hl�$X4j���\���c�$O��i�m��^zq{�<���5t��)��<>�XP�'���y|u��3&������+�����zKOA��K�a�eRɍ�*�����T>���a��i��a���K j��T8��z��I5�~a!���$E070���3���Ϯ���yk�v����I]�h��o{���50U
ңQ����z:d�2�Î�R��ڛU�-M���Z|F�Ý?���*�\?vA����q�}�[�ah�	�T���CF#�)T+Dw�f�)P-��PB��7Z`Ҹ"��P�
�4�.�F��k���:-�h@��_=��d�f:\;�\HS9�����=�h�����]�,�������� �*�!�rt����=���p�Q
��!���/�D��8�*��E7S��	T����A�9R�F �T� O��ϙ��o�j4�O�!HZA+џ/�#y��@���Ͳ\F�`�����GC:�3x�2_=�(��#c\����'�>��9ϫ�	5�h��^P�9�	���W�9���TO(*V�a?$C�܃�����ƧvV�[�X �Y�hU������"�������B/�9��{4`���!8
]��M�i���R������g	 ������G6(�g|��+KM?�Z��}�`/R��ė�q�T�GD��?��@�+�f��%��^�'��Ս���T?9H8"�H9m�7�3�O���`�%�Fm}u��
�2�ﶜ�~j�|:�8n��>���خ���&P��#���m�	�}�g�֬&6o����GJ�4wFB'nn�����"��٭�O���bS���� M�D�����k�ǣ�G�s���FM&^Ո�k"ʈ��΀f�a�Z���a\�Cgz�S�Q��[O�]0���\���b��[C)W��>�T72PZ�2d�N�î:��M���D ����D������E����I�9
�S�Y(ycN]c��?�<5(�Q��L�����_��Wgh�@-�#M,0�`u�� �'xD�Ʉj��6��Dz�N_��Ll�{%1.�	�L�}�pc�֭lt���v�7du�I��!�܅�R0M�Y�u'�9z� hG�U?���K}|j;��as�� !0S`��&5(�D�K�/�a�Bh��7溏��.���#P�,�E}��ʈ��|�&.L
S��9�&#�Wgi�V되
;�6PB	�Ùnx�m/ ���q�l��Z�$9x(�+	b�y����w�X���'���HQLg�}έ!���!��g_�E�������x].�eu�B�j�̧������8���H�$�5E��\E��:1y��,�!b"�����L�����ꐏLq��������ѽ�Ɲ��eљ۹f3�=�PBh+oz$�N����1M�*!����ٓ�':V�)3� #e[I0�������W$��:Q'I��&J�ІwYl_���3��q�R�L)�|�v
k1��/+D;;�V�]*�8q>獝����R���'Ӯ��J|���]�z��LI��Jezb�p���6�z�&���U�ě&D�c3��q�`9e�+��hin�N�J�Ի<�'�]ò�&=ЌT�t�uG��q�0�n�d.�"4Z	�͗|Mmv�c<c�v��ݯ��w��T��&�����훧1	�-5�a��}��?D�l�n!����r�^�� �*�B��2�T��^q��n�����_9�U��!nL\�ĳϯv���t�n�d�7HK�cF�^�0|�`�R�>�7t�,��Y&�o�ݮ�zԯoMA �t��X" {��0�
}bt��D�+PV�����A���,\Aa�O�M�_��g`�s���k��{;m�Q���h#m����A�#��[�Y��V�� j�A�����Q��ҝ�3�KV�:!L����6�?T�󄒨M��_�/'x_���}a���fE,��uN�Upð�G�oH��m!��}�f���Z?x�ճ��%)�����Z�����)��9��]�'ꗁ��i��7�/?��5�MGv�  ��Zb%cع�ڔ =��JT�kQQi���{�.9���[��|�f�nU�� ���<)�!���f5́�\��O �P1�0�v�� �w��S~���Y)��4�0�qS�υ@�J���^���PWbZkxl1꫅S�d'�U%%4A���]~����z���V�&�5k�@T����U�+����-�b�N(��"�I��i`o�O��Ա�+�+ل�$rD���R�c�(���U�@�"
I��߈����)[sS� �q�Q&t��&��{�8ᥗ �l$Q��5
a�Wv��x��Ƙd$� y��C!h�WoP��z��bd�Q������y+�|�Nw,���0hh���4v�Ʊ��I��5�t��u��;��Y�ꝺ3�՟�"�!)i{�X>+:3����ڦ�������v�ˌ:��g&�0�����s���h.��8�8�� =�Ԋ+~��}?�BI����A��ԃ���R��4�T;��gǗ�x���B#�Z�x�ɑE	Ux2�C���_l��@��s*��x��\}{t�����gL��dF��9-�l\4#�0�����\����\x'$JQB!xd��k'(�����*7ǿR��T�t��C�-���b,J�*�����8=���H)ޣ���.�!�����	��<`��c�=xTm�ipɼR�2Ș'HoqJ7���Y��f��s�aF���c��9��r\"����H�qm씞ki��.�k�!�O۩f���7*��V��z*v��F��d_��$H좩)����hVu8�J�i�Ub�q?��.,,���6O8�`��Zhv���7�-]VjzbU��Of�'mK�Õ8<�z��Wp�Ӗ���\돞y�Ob-ܽ�GW!O:~5��Ӻ��ĨpvDF�聑��}�M�ϝ9�aO4[��f&'\� p�Z��*��`��,?�����˷�<�),;k%��#�h�? 
?��Ӕ��?IL����ܮ� ��S�f���轛^�$�Y���}4��yKjR��M��i m��1�NP�L�T6��(�̰�6W}����vU�YD��]�H�3��n��f�
"/ăcu��� �<-�xTt�V3/"��
Z��Ϸ�a�hI�C������LrZ��ւ���8�h�c׉�7�X�A�;���{\�˺F���>�ȶKPqQܑ>/�}35zSt�@'�IT<��lL�h6�		*�DL��6L����tb�P�����j>X�o����3�՘�s��%��=�A�V�lEAQX �w:�Uk:U�\բ���o��An]SK1S���x-��L[�m���1��`�&A/�<S�C��Z�;�<�����`gc���k��Zx`���s�D�v�BJ����}�0Qĥ�����2j
��j
a�>�X��JD���d�51�g�7��k�GK-��l~����va}����6�L���
ό��
������	����"����9�V��Y��RZΈf���-oR�
>�Ѻ��o�4��4A)�L��r���)�\�W������=Km�ю(�Λ��h���	0��Ã�܊͹/�E�c�����\�