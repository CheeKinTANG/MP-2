XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v�����ySb����cug����/4�6Q�v�C�H�{�TH��l�0UoIa I%��qN��h�M�5��j/[E�h��A7���3�E�l�?�7��{<������Úe%.�����fu��9�Kݑ	=C��[%Hc�@�/޲.sA�i�m#�2ݖ4c� 4��  +fڅ�CͲ�k�7��D�6�!pU�b�B��R(�m�����)�h;�*�ɯ���ٴ>Ԭ�p#u!@R��h�Ҽp��R{�᯸G�� �O�ב�dd�����(���U�k�O̟��v/�������}N��_����%�C`"�m�ִ�r��o���\��+9�`Slc�)զ�ǃ_Q����/!��ym ��G]�rk��9I�2;���8�w�E$m��ӫ�UM�y��t#0ӕ��Wb5P�G�R���)�u.�Ԍ���N���\c�#S�G�M���KG��5@bǜ��R�����s��j��m[+~Z�������[-��W��#��GV%��a���OJ�GV{q���V�S�L,�O���V=j�}��
}�(�Zk�اc&�D��yb�>E
��͆`�~��'"P���%.[m:4��=&>_c��j��ٓ�h��&��<Qw�_t���4��H���$�!�}Y�k�h|�#��"���kD{���@Y����]��`$����>��,Pgˈ&�v��o\��c9@<j�B�C�h����k������aЈ�k�2�r]h��IdP?�lA��mc��.x�.� I�3�=9XlxVHYEB    da59    2e30���)�C�be_�a�؉~��Gtb����A��4�;�אD�g�47H�x�~Ɍ����"Ȭ���)i�������kD�RG?�D�l�
s���_S>�>����YR_��¯�LE]>k�6�	P:g6�&�������'���j�I��5Pʇ�O`R��ܼ��9"��p�e�z3υ���H�6/>M������ګ_���7��㑨��_w[m�P�F<���QJ:ux����G��T�k�)#�
��z/����D����6)ゃY�Z}�l�|�_\k�n�ڢ�LC�U{$]^�ͅ��F�T�/�����*���ܮ��U��T���x���l}7/x�0)�����V �S��X������}i�"�.p?j��(�T�Û�ٛQ�G~�>�zX)T|�����|R,X�yd?a��V|���.����IF��d��M��"��:W��7��#�VŪ�P�M��}�kq�����)�����6��G�u�a���fj�U��+b�Ui�������_5�o�����u��,�1���D������y�x�~���C���(�~܁Q�lã.M�����,j�\�����$"�.������ ��Nv̥��9�zGM��=i7�����tי���	���a��˴�G�Y �Uߩ(�P2:�fPsD��Y��OL^��\٤�M��»��#SrH��酒�H�r�C0�kW����t�-�k{���?�}j�&Mz�Wa��U���!^>EK�j	�FuϷX����"k┮m���o�[�� �����Gf'�dO�%z�@%�^����v�ynfן��&Z�C��:zx!gpH4(�
qF2.R�WD��0��V�G\Sr=��=��Q59zR�����h3 )��Ǎ�����ȼA�DQ���-���/U4�
ك(�2�6�9D��oB���#֑X�^r�T���$�5��a��X�~N�-ϳZ2��1�<"U82MZ8{�b�b�j�Y����!$��
�_�g�|���ÿ���C�V���v5�k��� "Uq�!׺����CǶ��h
n<}�����Q�H�
��|Cu,*n+؄�5��d�J�J�.�����'X�J=��nkl�����e+�!�3����T����U��p���#�bl�t�)�,��b-U�V�y��{pn����-s���ɵ������X�4%:򒼌y��Ilo��d�2nL�kJh}_�rsS� ���@�k��@��q_37	B)翣#�NG�j��:-G���6����K������W� �s2��̔�����M]�>T�4i�g�F�����7D�N�Il30�C��$Vh?�r��3���v��+���J'Ү��hQy����VEu8�p#:�����\j ����?8G�g/�o��@r�����Y9��X��U�r"p�v�.�|�8��q�5��������93��"��G�*�(-�c�?�j��uh	����i�)�
�AHj�����AY���M����+�I"��Y�F�R��J,�yFZ�>��K|R�F�q���Ǣ���^G�|�
(v�⼓,B�R�nY�������t�Y��o���1%[�v�XB��h<Z�	���;�;�`�|�q��<��f�(C��M������s(Yn�ɭ\t�Oh<�v�51��[��c�0���oN�����%Ƴ��66)YX7��(�n���d�	Co"�C[$zI�R��r~իD������#?{���ѯ��2��'��K�Y:���.��-���i\8�Z!Y]��K�!j����7wZ�SG9-b׸9�Y;����F6^Rb��)�@E�bn�ͩ�C��Ŕ�����"Ȣ��;�k���|X�+�׽6�W��0�6?�HF��{q�j˅D�<��h�P3���[SB_&��Z�Xg��`�w��$�^�c"��(Ǩ�Bs9���i����4qk���.{�Zu%䃉Ӯ�o7���C�����(�9��}�ڂ��ؓ�P#�>����4����;BJo�>�5	�49���o?g��2��X7p0��?~_P����ސc��x�L���,r]��*鎈o
�v���}^�t�q�F�w�c�%Z)��3)�5:&7W�]j�;P�W¨S,���6��
-K�3�$�&���2M�](#�N��ې=�-:�H��
�	j������ָ:��H��E?'����K��M��쑤�����%Y�O/z�ms��pV�"��8�yo<��3��*z��ӱ}����j)�q��[0��Z56��9¸s��L1�i�cl	��[�hv�L��<�4��:V����|d%	w
n����p����g���]��-�������Aq5���$5�o���U�Eq�qu%�|�F�{�?�Z�K�����t���ڦ��٨~��ب#D�@xp�S�J�Cݔ{�ab�tM��[li;���@�)yu>Ӟ3�6�R4Ȗm���[ۻ��3�f��xS|;ZB��Qh٨�;H���B�����"��cY��;��3��%�<�ԋ���N\��R�\�%��:��F�{�����O�y�b�]=���8@
��Fg��a躪��8[v��` �kA1�+��pjL�S,��.�|ٟ�F�gw,�t��HՎݚ��<Z�}cS*d�zn���n��70��>����Vn{�3}g{��`:�+q(���(�4U3-��5��ܔ̘b���b�W��F3{�� ְ ��?i��?�:�MC&��[���N�مvE���D��5i�0�-EE�%Ƨ�A��X��.�Q8[¼������ �^Rʗ���K.m<0���~���������v=R5�U���gZ�t#2�jMM�!���鸈Y;2m�� �-��K��$dB�7�}̂v��:�S6StDDWY��v��X�h��#�A��ԥ���lLh	��zAQ�����e>�!�kg��]�Y	��e��nW��PUR0 ��1�J��C��oP���{	�j<��`�˪�Q���Gq����d�m�GC��ɝQT/�BI��0V���b�*rd��	qcَy�R4�F��ގLd֢h���-��=x���(�OﲊJr]j�~Y�V4�	�����T�)�㬨��Y��Dm%/#aQ�I�@���O;� �'	��[x��Q/v���(_#F��e��2�]ZS��j�>~%�������Z��Ŧ��$���o�PR�*.����*;3]b�'g����~�P>���B�1��T�l�j����ʜr,6���D�9��r�����O��o���.�j��W��Y�{A] ��Vt��j+,�=�hhX��6e�#L�S�)���O��m�8��_�=s�	d�������D��N�X�2�͢�|0�Ft�#0�`�X�N�ɫ(\~W���9�NrC�J��思X��}e<ZÁ�h�hۀGXf�T��Ε��20/�ԃN,�s��;-�9�1�R���Z��F�P���K�扰#� ����h~�����R���+�D{���U;���6�%"L��Č���L8���ۈ�Hۉ�"EL��6�T�E����s����eK)�/7��nߛJ��9�����:��3�e�✙ 猦��1�\�����$z�QG�@��b7������yd�\�m�;o�)-)�=T��� �A�Fb������ X�Y��� B�s�]����Y|4"���^/�X�Vt��z ���"v\����[ԏ��ץ��I &�FhtM\���6P4��V�kTO(���$��k�5�4���CK�D/�j+�X0kW�1���E��ze~�G�&��'i~֪ �7���X�V�H��/Zb`�>�?4��8�' �h������48Y�ӕ!�6�����f�-�+����4�����`!po����o�L�,����TUU�[B���"���4�D�Z���t���Q����E�xV���(�[�ʽ��Ζ�yh��S�˜�iH���іmV��b7a�K�6��@�"�̦)���S4'$�U�m������r˦%�]�����J�C��	�1�����^ž/q;-�n���������z�U7��%֡)��c u�W��4�O1��?g6���6 ?ȟ7�w�b�N3� G�5`ujf��^v��l��F��Sgף��/������Z.�AW���<o������;D��Bν·�� tΒ���qo%����dj�F!d�+�5\���ѾT����ӀR�$[K^S�=�Ĵ
):Ð+��.{@t"�����zQ���B�;A j���N�R}$)� P}]3~u�)<*��<��2MwY�C�'���9ЌrWҫR�(p��4v�r��F��o����z�ձ�;�ԉ�PJ�PD�:6
'д�B����6���x`��47\�̣L> Іy�-R�̹X�ӗ����-���A�}���ˬ˜�r02�J��������|:b�#Ѥ�]���&ɛր��h�`ʃj�Hɜ�Ո>8+M��t� *D�*�?�H��_��v)��!ɀ?��L���6ʑcn�_�/Vԫ��ݥE�ndЃ�C	�+~�22��5m���� ד�9�+KS%M~ߏʀP�~�Y�H(N ���>A賓ʤ��ۀ�E½�hA�n=�a?���@%�`i�}��_e��u%.�Ϟ�LSi<��rg���d��_O���.U�V���@;?�L,H/�%P௾���^��F��]��v7��P��U1���Dr{#���z�ه�����5�G~���� R�	d�S¤p�R8w:��"��I�cկB�śMfQ�/�z\y�t�̝�����Q��66�Z@W+7�ؘM�w�����G
%=b��m���h��������91���ᶖ4Lc5������kՆEZv��Hy;���.���X��q?�7u����+�g�����-/����+FP'B��V�N��� w��D�	�d�_�� ,L�kKXL�
qKL��[,Xy�>yGN- Uj����:t�Y� �an��8���y`N� �j����̱0б�G�^Y?/q�X��߱�֋љ�Y��+'���������8?����jM�]�m��� ����>F�eA��d�/`��:མ�G�I8���w��=�:]14Jv�?�c$���I��Qvs6��G�H��v�漐��[i���&R;��L�6��hIێ,7me����^9"䄸�9��oB-Lr��,�RV��+$�N�c�XO�֊�t�ƽ�.�Of���1��X*.���� _���<G�8��B2Iΐ��k�C.qQ'��]�ƐW �O}t�"�����n�:<gŬ)������F`<��]�H杯�Q@��3ʌ?)rר���-}�a>��!��h=�͵�3���)��)0v}�i���n[���$"�1��O��g�>���z{I�NZNG5�z�H|"���;�n>��ý��5@�v.O��x\0%U zV��B��Fh+���0��~���idj�[Q]T��U)NgS�lx�_E�PKH�_�v�����ΐ��5�Qό2��~�Ɔ����Oq��C�us��F~�Յ@�×�^L��Ƒ~�;�+YZ�#Y	n;�:�$�ޣ�Ć��� ��-�wTW*08�?��0BV����6��VM�Ą��@�)���i���=�C%��ύ�YE��-���0��ҷZ�<��:������5"��WK����cp좥���f'�g�V�.	r{����Sd�m�1���+���,4)���L��8��p0{��ps�zט ��8��7�G
�B�ٸ�g�]��=��Y�2>!P&�#<�pP���z���������~�ݴ�(O2
� Vd��J((Ri��A��}EF:/�ej�z�X�����^���[*���	M�z���~@_�H���,~�K�`&5d|=P��L'Xx��F������
����;@³��J�xy�Qv���EiG�'�R��/���=�rf��^���}@e�-G���#�K8LA��$��F�\?����O!�6Ї({L�lgl�¹i��{��[�/k?����	���O����SյՔdN���jmd��?q��8���!.��qX����*��c,��P}�x���mK��FtT��J^�G(��~��c%�$�Y� ��M��K�Y�2�0�R\�b@�4����-�7��z�-7s��]�s<�d�w�\�؈g_{�]m�F(�~�;r�
 ?��L�2��B41Gi�\�.b<�ܨ�>}�ƒp����Z���Қ�B�Q묻��^ a`zS�/u�A&ɯ�e��q>v�͋��e� ק)���0��((���Qb��O��{���*^qX}T.�l��x]D#k�m��k%��e	��,&jً�"��>�Ւ5Q��ʝₕ��:P��/�m~]ЧZ���3��=E'�}�)�!�"X��`vf������Rw�]��' ɘ%p�Yxi���/��и�É�d�3�	#\)�����b�wh��W����Ĵu�IJ���#�1)�J�u~���:�g,�J���5;����^?xd,�I(����~:o�W�;].����Sz�>��G�/A�R
�0�`]��ʆ�X�K#��Yw�����m	�jp`���p�#(RN�՚����u0yk�}]�}T����eb63�3J�Kv���-b�Jj����%����b��B^V��2�J�s,7������9��g�ʬ�F�$��hA�cY�_@*�dZ��p�R��(G�	�Nvq[�k�����R{��=���T�HQvK��F��|���*�5�f��Y�D�"�馆q���D�<�w��f(�UH�$[x=�ہ�	�k�'��?�Np����:H���8���/&5�-�*u�A�h���3���r��?�N��pA����=�������;��]/��$�HRo꿫�}W{��#Ұw���r�̋�2�lK�߳�MI���<4���>��N���#!b�r���5��vW�j��uN�\%IR��kJ�da��^lK���d��l�/0�x��Oy�+m���!�:A��V�F��+$���dt�#4X5���������K���v�3`SH��gڇm���a}:`Q-|��1�Y\�#'zN�0�z���M�Ƀl��N.���tͰW�)������7L�{LY~8G)�"M�>Sgo̐I�ୀ�`L����$�wLA:���Jf���*ӽ�6�_*J���r�E!n�P�Ɔ�j�E��N���Ǩ��\���)�����(ei��'�p��@��9�$�U6!=�Ӆc~z(����9|�T����"�e!��.P�z��~%]����A���2���8�%�������.I)�Y?����O̰yE������G�-ya��J)�sE��p����h����8��3��kı��^x�cL^|�r	�"l�]�=X�_^.]�M2�<,&r�X�,�{dxn�^�E~3u�U0���뺼�79�~J/0:���,�߈�蟎n�,{>�q��xf����E����qa�&�p����(�&��=�Q7�\����9c:��y2�x��ݝ�EM���q	y�u�M��G���fy룕u���֪{g\)���_��5�2�d�;�s��[k��кBͰ(��2�p�@��u	����: ��e%(�!�GO<�_���!eh\"B5��XSN����t�<���4E��KY�+�Q��b�O-� ���K�͒��7�y�s^y�Űz���|��M���Y��寽�ǚ���_�I�{p��w�#���@�0��l���A�!��؛�I�ƚ��r���BOiY�ɺ�M�=�}r�C0��ϴй8�=����~]Է�����;�٩��v�/���82cY�n��u��J&���?�]z*��S|@W���3�"39�zv،I�Dz:�:!O��h��k3!<}za�p��Γ�IN�h{��>�S�<�C ���G���쵃�kN!~̹�6�M�J�΢��4��{8S�5M|̙Ǹ�(���Iy�I��S�$��s�h����"�U�I�;@IH����5�n#��V5��S&o�D�r�Y-�r:�hg�+��!2	ͩI&ؙ�?N:x/�X�ln1ͭ��Q ���QU��"��Y3k��c��]2���'X&��j�?� �B�lK�i� ��C�m��	�?*�cf0��(]�@")�,�v�>����q�b�����(�QS���.����C�J��%�8C��q�f���� :���ċ���W�I)�.���n��k�,�ݡ؛�4�HSk�[����j=�W��3V`� E*�6���b3Ǜa�«﬛��r��Ty^�.L˚$w2C�!3�W*�Vm�R��q�Яp���=}�Յ��@�����Y�5�390�u��O&��m��dQ>��C��僺TB�;���d�V�ՇbI�0�q4�q_�>W����2�,���SX�/(إ�=�eOw�9���E�G��m�'?���msLI.�\��hIO;��1�w�/鷿���_Q�pZ���a󋡊�Uh�U�k��KY�Ь!�a�Cpa�("�5���=˜�~���$���H^#-9P72�~���P�(Vhzit�]�����h��N�] uOH�w_(rg���U�<#�R���>�C���8����3��5�1&��7#��8�ж2��zS�d}��N҉W�F�#�?:G�R�p��YO��b񐹬C���߲���
��:�05��>�+�+&��mT���Gs�j�ESQJ����E4-�`!b�����?g�|�"*����a��
�S+2��Amx��z$� (�Y<�#	��P��+G�x//"��̚��.S�[[�n���
G��~��w�_�9*�50Q���ri�flw�D�%��V��F�ˡxv�+c)z���АPy8����N ��1�s�xZ{K��#�����t#z9�3YnK���$��;;l�P�?:`�#I+A�j��g��.b��~ M;���ӭU�]/�)�X�dc�����T(��V�ը
�BA,x-B�d��?����}��~W�
�G��mu=-��L�����9�!�XeSl�$�L:���qʣ{ͷԨ�T#���QO�����D��+z}P���"�'%)���8D-��wl(�9�$*�q���}Ю�N�Z�{_G���s�>��<{D:�䱅���� �+��FP�2)�u��FM(��B�wT�׽����H%�k�o���?�B�f�AN�?�&�̧�����Q�܎����G���3�4̈́P�����E��O�(�y�Ǻ�@��yȪP��Y^UYf�-��G���?�9�2c�үy����呛�ȣ��[�`ru��l��Ǯp�M�v����j�w&��5�h7�S��3c�'���!L��k�
8�E.`����P�m��(�U���?w�	�谼p�֧*�������3������0�e�_o�Mq�� ��R���UA�oL�U�����}�)�����W�� �65�Ϟ+�mn���oЅ{/vo�i�?'�z3�}9�L,Bny�~�0�r��t����+Ԧ\zG��i���#d<��
ɗ/�y$�c,t?��Ҧ���۽����U���8N#[��D/wm�g��N���<I8�
����8Pʿ�Y����Pp���["|�"�HM�`ޕ��*�4�֌�����}��	մli�[Nx��@�]�� 1�+��Ր�zN�QB��~d q�A�5�H闒YSJ@���,���Y�azq�k���4��'�p�vcC��o�JR�)]�7+��U9	�����:�Y
M��r4Ʃr��l��L�i�7l��O;P�O�:�Ac���ҝ��5i�|�L$Fw@8���[2��t�X�P�����QL�?΂6.��R��S�G���������Ԓ��1��ݙ���.��bܣ}G�?���>b���8�H8 �m�oc��*��Aq���su2��OP�z��2,�n�����y6�r�6T8z�Y�p���\C��@�߳mI�[��O���"���՛�-���Yod���RW���x�����I�4"ߜ��b&;��⍇���v%��Y(���+K��(�C'�Ne#Pq�2�k4�z�|�ZT�HP�a���U��:�"|�L�>�������S&��)&�8T�;�C�9���
��#Ksė}�'�Ǟ��EM	OX�B)�5?��e}������e�kX�sf[(����G��*��RO�&��[՚)��3�/��G����e��B�&��S�ň]X��[���Z���*գ��H�
zL�QkbW����� D�؜��w�U���������=��[�� Lx�b�=Fᱜ�2�c3?i�L��h�D�%�M��־�F�G)z>r��ۥM["qU[A�����5ɝ/y
���_�9c�FK����'h,�\�	^��$�4KS;0�d��*�W��ӥB}��a��.,޼D��,���ADW�-L�3�_���o��5r��݄�����*�Y$/���U��KN ��1-��P|I��Ҟ�}�q��,ZYS��/s�C�j�T�Y�IDR��ų�=]
��Q�
��-�8���ڿqEϽd+^	��i�K����{\i\OI��F�������\UPQ��[����!N�9tZ���*گY���a��z�V)��6�gI�(�%�p.�$�z��/�����ofx|O�?1�f�;s�K+�!�����i�cz��6�>Z��������=VF@%�#�ʧ��s��תL��6���k�A\.0���Լ��i���g�Q�\,8�F�Q!�
� �ui'�B��9nw5�z���N�@���?'Dv(Y��2�d�FO(~�[�z��~~ϧ�^�Tu��Tc
�u��p��<���u��\���_�)��2�݉�h�/�Xx����6����&Q 8���!�iZiA�����U�z��fOx���ԯ1Y��eX;!z5�IPf�)�Ṗ�eԆK�
�?*�]���󰄎�.� ���ie���OJ,��cƉٮ�D*k�M�#��n`Q@��]�����	E�'F3R������u�|�kfK`����!����*	���S�	;���(���E`�ж%��ʞ��Q���	����FS (j<���L_�r៼V���kكȀA�^
���� ����!S��O�r��M��('�:ȳ7��jş����0��䡃u,prj%�K�T��3�ѷ��>(%��;�;�"���ޅ�bh�G�Kg�z���)V��B����d�k�߫C��f��W�q5��{ZUh�0G���p��#Z�ԓ�Δ�J��:=��%sj�>�-zai�$^L�c��߻[�Ӝ&���æ��`n����1�z_��֋��X��6���Y�o�!-�=�`���z,�����8���L]��T�����	*��b�EE���{�y�booG��*xi_��q_J��o
��ऍu��8�{���w+��I\k	��1c[7�}�w���%O�<Fc�XD+;��!h�1E/�55a��V���o(��q�����e'���r�u�{"� �	@Θ�ǯe<+�QӺ�`}K;Zu�~��ŞX�O��8��$���ĺ�Z�^�|ai/W�#�8�i^a�F�ր�m2��4�8+\