XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q`V�]�mdɶ��R_��n�ґ�Ձ:�/��K�Q�Jxc���[η'����m���ap�ư�C�6�Xi�:�-��﶐D�5s����~��j1�y$Gn�I=����lԷ�؊ӡ��D��f.�� Np +�܄V"��4��{��̀S=�[}�g���B�s~6�xݯ�.�kU�,��J���d��!�<\ρ�%ۇ�!Ȋ��W�2lCS7%�>|*��k̠>�����{VK�,��R����l�?liW4V*>�>��6���p��L?�G*��E3������~�G���?��~tg2�e6U��;�������*�6����i�����E�J&ɛ��w塳)fCh�()˜7�b���*���Z���� �*� g���P-�C_�u�w\w��~`l��Nc�E���>��/��h�\��y�����5?�pJ`�k~'ېFt�V:P��$������|��P!d�D�&�h�.�)sc�Ҵ{�����ʰ?�}�'w�P+� ����I�a_!c�fM<�o�w����S�p<�&?p�����sS��קꞞ>��*Q��qh$�<B�d@2j:C;p7=���h���a�e���asʘ�)���Ge�mJP�O�˭���Q�+�%��0�b}50Ɨ!���8L�O��|�P�=��
A�*){��	�� �B�3�������H ܮ%�ʑ�ң��L"�.� �d�?H���,���O�!EL����ށ�*o<a�˰�)2��홊XlxVHYEB    39de    1170,����#������z�<�ML���=��&�<>�;��>ۣ.,��/�8�]W͍z���&��~�ƻ�7�+�R����>%$?Ŷ��W�4^M���W(��֨b���b��x��{V<��A�S\�dz���YC�Kh�zT����鄏��fQF��	ǐ~$5�r>�NO����#n���M;���h��#RW�ɔ��N����q�o���#8c_�^�Y}׀�-��^��w�lδ�S�\�ݚ�>Vli�L�����~��m�8��m�r-x����&��%& ���AoJ���(bL�����*���c�'�ua3�"u�]s�Ԯ��#�p��8��V���5F�.՝� W�?#ka���!dO���Aϕ_������B�DT�������lk&�D��a6��_C!5}�&�,>�ns�KS2���
�߿Aٹ_��A7���v=��^[~D�1��s�:Y��:{�<�+�����aA�kul�&�3�Y�*�g��ځ` ���R��#�e4����х����pd`վgB6�<��G<"���� 3��v$"����� ��[��;�? :Y��rE*�5�z�Խ�u���6ppƣ<���I�{�|+�fu��]W��_N���q����M�f�ヰP��P�t*�����pʥp7��ox@�~����@��Eӝ
�@'r�>b�E���}Y� ��1s��⽷?G�K�
q#D-Ym�N��|F�ä�||R
~3G�#�E���Q%��n���X�X��N�%�M�)�����j�x3�7}�r�q]({�Xk(�>�^��y��TH�`��ݛjɦ�E�{�T�s*f@ޝ�������v���J}�~�{e�X�D�&�U����P`��%�+|^�|�wFT8���Vn0��1v����bU§��e/�	$;�����Օ����Ab��d���{=��x��`pI��1�n�7����0�N�����G'}~p�W��U��>�1Ze��� _+��r��7� @���+���	(WD�-�� ���=br[]�&��p�&b���D���yTE:�K���-P��.~�1�W1��{�S�Q�G��I��I3��T�������	,�a�ڨr0b×�Vԉ��|���T��P����Fe��0`�3-�s"�XZ�C^���U�y�M��E�Y'�����#1�և�E�!辕��?�i�ux�ե���p�قc�-�"g0�d3邥\�N%Qc�I�+6.���&2���	ß�_���Q��H,��K6�,�����T��mȥ��{~��:�&�����X�#@����ظ���l�)��a+ӹ���\iUVm�:�ҎG�x��]�ۂ� ��*�9�T[
.�C0���Hw�D�T�,�?|2�bd��x19#��p�ryČ�!������n� ����!�(�ƞ+��i�ж���=�c�qgZ~��2�[��X���D�k��h^�ֹD�RyD����ttM���y�h���w�C���2�=�c��R<�o�?%ţ&�\֐��O+�E��<��u�m
�c� �鑮F��u,����K�3~!c͌!�+�E2Y˱�yY��$������1P@���3�L� �*�������' (�Ђ��TK !EFtX}��z�j7�ȱ��������T�h�FW,�Y��[ѵ��G��wY8t�e�+PW�V�8�R�l�l�duf��pq�#��V��i��7��?y��-�Sr�+��Z�����;!"�C�	Ǟ6.�9�݈�:̩"b�2�W�;qg���2�3������e�ͨ��Z��,��;�in����bғ�F!���m�W"�:R��0�o��-Ŋ��$|Q��6*��&�ߟ��´���Ǹ�o�C���j�Ѫh���Uw�T���h⛹��C8����ܳ�J���zb�զw�Ⱥ��M"����5�k&��T��Ư�Y�)�)߇dI�A:1��~�C�A���S���'�B.;��V��m���@��d΍Q�M�6�ᩃ����1���ຎ)/%ݿ�����%1n�ޓ��}�h/�\9n��������"�ލ��t'WP�N�M�4�I�SY-ch�a�l��?�D&hX�&��� �8�&]a�d�[�j?
h�3���שyjb{�ʧ8K(L����`<{�(R�y�a���̿�Ī����y���C�T�M �Rp���� ���q�i!�K-Ao-/C�3��~��/�BV��h��U)j�W�S��an(�HZp�a(��Zή��e�G��HC~��A5cEq�ڠ 
\"�v}�P���t<T=�q��5����D$�t�a6�Jh{��!K�bُ�o��	��h�^�._�D��<�cB�XRѤe��2]�S�{\	H1ˢ�3ݨ�(��� �'w���v ��x�����l/��+H(P*y�a&1��1}��uR.���o:>�h�E<{
��$��J�7��e,��_��U��'Ze�z�e�_��fɏ<A�1O�GH�ݲ���{�ʓ��ጽ���o���D��5���I/ʱ�<eɜ�ꇭ*Lt��L�7���Ժ�ڀ;G3��Ȇ	�[��X}�/u��	A4�ǀ�[/wxW:��x����U���\8{��c�T�.=���9���5����۠.�sr�px%`*��g9�_(�	v��1�]��u����˲_��㦧�Z�
ǖj΀�~/�n���� ��l�o�̝��Xs!|�~�PV͕���OFʋ��F���)�<�gV�g��bF�C@�GC_rf��r.Q!lO@�V_�E���k[��I*�{K�_e᤺ |,EE�� �9JF=5�ZA!½Q@U�i�HZ:J���:MQS�B�!���_w��ձ;�]��>tc4�
�꾿C�5?wk;�Ѕ�;+��ywđ�(R2s.�2��u{@�!��:���s��ac>�~=z/y����g8D��R�9W��PX<����ް**�u��z�g�)B���a0�?Q������DkN��WwN�����/�9�Cz�ۖD�K4QqZ�u_�;�W��{���&��␩0q�Nޯ(�#�]�6Y �Z+�R����ﲴc&�%���U[i��V̚�{x�|����a$�e���Dtz�H*ez���E�o*E{���UATd:�M_��QlL:��h��+�0%\rOEz !�iN�.��%�"�T���v�o/���^�=ި�Ȍq;�	������c(�T��&�E�tޏQ}��������M��h�����;e� y�H�!wq&���Ro��r��+�s39�6�ap����6z$J*ؙ	sjg�XP�� >yᡁ;/�\jH��m5}2?�V}P�]���G�W\^r�uܑ|��l��J�g�q�)}��ŀƶ�`w��ĩ�V5�P�괜.�yJ���W'l�T����z=&G���Dk�#B�'�M`e(���들������*Y�%G��l�[����,iNh�-�����%������spJ҅�j��9�O��o�	�Z�k]�X@)d޿����]lyK���%�9x� � T,k���ٞ(�H|&�( /��Ȁ>��������i3V��Zگ��D%i%[IIe�
8��ԃ�d�]�N^�^�R�*� 4&�!��L�3�»-���|��p��?1�L�=q|�Fَo�(�D��TȽe
�Q]P�0�ߚ��[�w��O���S��O>L4���廥6��&lR�Aܖ�N��y8U�����G�>ؽ�6~�B�W���M�R]S�c��V���}�}�hC��kLua�D���\t�����W �;HK=�����z�镦Jt��� ���IR��������#ՄuVEǠJi�֊nZ��dkh���,,�@H-�zB�$��V�u���N��e鷺P�����%�RR�9�/�?z7����:�X%c�<H�io����Y�b��*��������o�}��&���ܸ����A���$�Ь��Y��	�ʞM�S"���Yz8
��l����8��D���J�I�yN؋J�E��I�6��;�,��KP��@�g�դ��4��ˮ���/��g��m�@�*����	h�u��?BH�S���5�mD���
l��R��IjGI������LF���X%q&Ǆ��ie�^�����������ץ{���0�E���Fp���"���M��%�M�*:"m���E�
��q���sw�2��!Ƒ'6&�����ɅzGt�5��;R�8mITԐDO�cwQ��3K�=M�y�@F*<�F@����깼8�� ��uu���e�K��7��>�gʁZOd�Nb�WC�E�0�膏���w��qއDk�Xnw���(��4�����Q��!��T�794