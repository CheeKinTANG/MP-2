XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I���*������/
��q��&"�{!E)N���AJ�m<)Wx�6'��$ۣk���?�P+����_�ǈ�L���5�oV8�2
�`�'������Q ����]螾�UE���A�_�s�V�$\�VJw@n��P
�L���ĥI���+y
�ʱ���x��O)���Fi��#g�����z_�B6�1(��i�VCC���jx0V�gH7g(qʂ���o�e�,rEv�?%0�rƥ'9i�f�\����l'lN�}�}�췛,s�K�3�2d��GnS�$-g��ѽ�3�CJ�����v�i{�z
�2A^����N����Z0�6���:<1(ƊH�
2�GV�֤6�����Ѣ��E_�t`���`Κ���,��FM�����7�k���ܮl���õ�C�)S����t�Zx���(���a2u欦���ޥXMt���l��ȁ/��:O�O���{��j�A���'�,��v�z��z�eo�"�_��2-}�J����S�C��x�[��������-��%CRu@���`3-c��(��'ݍ� l������S��P}����q�Nu�p>?�VQ$�~	���G���Z��$ -�����-\S"ZK�,���;�O�3[`Z��q��{K�X�Ĕ?��P:�Omɿ�b{�r�&�){�]��Bj� I4o�Y�+�����M�z��t�B!�a��Jre<�Ɇ��m��Xk6�AJ�w�������:A�H�4p7tm@
*��nJ�XlxVHYEB    5224    1740^t$���z�c��N�%�������%o��F���^�s]���1`�w:k���0\�$��J��|t�]��[Y�Ǉ:Š��"%��29�V�};�>�D����c����ʶZ3��B	�6��Gմ��OL��i_�v���?��#��)"����e�xK���h�tLa�H���4��'���]�)7�/\5r���tܑl�ī��[��]{�Cn�������E���
s�,_7� N�&xr���:"��� ��Κ��7)�י �bͷSU&���a<�0�2�w ���2-�?~�dz��%�o��uN��<��b">VhTZ�h)�k�<�@�z9��%��c
PC�v�f�73���F0��B�}�������p3Ύ����u����a4�C�ҞzW�+=Y V0���ZW�fW���5Y�Z������VuIY���]}̓�1J8Y\�EKج���"�؞�>��dDiw�	PQtQ)b���b��r≅�1EL� e+ }��-&���4������27�f*����Y91����+=%�-��id,�U{�@�ũ|�uLE�1f���<��a�UL%�f�W3�4TҎn^R�'?+��a����\�&3U~r�G�U��En�mW�ԇ�Mp�D'2�.�5YfΜQ蚲:�!�}���r��+x��F�3�W�3�o�G�$������n ��>�IɆ��\�/&�%͏�-���B�/�]�<�<��ӯ&U�qM��F��y��hd�	�|@{�"�4�F�r�^�WoC�3t�V��!�dL��jP�e�oA�Y�ԉC
��!yF�Z��)�wv3�[�NCOk��Va���YU^���|�.���x�7��Ɉ��E�R>���%��E���1&�W��"�|P��(޾�ྑm/�x�7�r��?������IK� ��l-��M��\tnL$����g�19��X�!��Lw��Wu]u�,@�YK3�M���	�Ͱ���T�К��MT�q-h�5�gH߁��t���n��N�뛦�u�fۑC=�&��D= �f��=���sc����Į��e�l��I�3�i1n�w/�FP,��F��Jy�w*i�%���(�x���8K�=�^]'��V�R�7O�3d�h���g�����]e�����S1�p����d�UqW�\���&!��q��1,�׎DN��"Í��r�>%��b�oF�F
�5��R��!U;�#�Ǯ����L_x:�C�:
�ڗӱs*�.��><�|M��hz�2��#�ǋuH��f��l�H�b/��S�_"̯v@��М�QR� ���&�k�c��4����5	�n�p��Ts�Q.��������X��j_�Gd~���+�<|�Q��<�F�06k��[({?>K���A�������IK�i��pV�����Rc�d੡0��zU;�8�RF����Ԓ���ї�ZJE�c�Ĉ�(V{�J�C�4���F ��E��s�H����o��\���3��
r�����Y��h-ep�s�����Ɠx��=0�k���l��S�gsQ���J;�llT���{R����(�5��-s��%�w�>�v����e�je���I9�,J7��|�<L:8�at 1�~�yǳ;��Qw�W�򲷉)�ΚuW�~2D0TX;dy��Qf�Se��(�-��/u�{���v|�q�S[|�+�|�>���=&@�}Z�Q��Gp��BC	;�uz�0�eN����Vn#�d���ϱ<�>�J�bnGcY}������n;H�|w+�7~��m��AwNG��~�!J�uo�TJ���₠u�f�xY���N�d�I�z�z6X��%�Bs��u���B�PY�r  Ƿ����@��p�� \�ǐ�f3�t��S1;+�<���og��ڕ��D�P}�K�:�x�|�4�gGMD�";ܑ��i}� �>t^���j�Kt��hh8���pW���y�"�{�z���um�SP�8T�o;����
�$k`��q�xC�7�Z�i��5{�6ep�q�-��
�(F��a&�"z{A܀.,�Ʉ�I���]����7��[x�ڋ-fT�^�T�+Y��]N��:�"�u6j�X+�7Z�)e��ʔ٢Bp��b���Nܻ��f�����yY�W3+��8\�����;�1�f��nԩ��8ꅳ����O�R��лA���Wu�2�0�M�N9p�����J-~i��UJ}eB�\oz�.uFş�Ź�v6��r7|�C�U����Sҝõ�3���t�do6u�����1o�U�[\��x�_=��d���h${�;�C~��IT���%�Bv/��`����F�M�T\B���xب�ܟU-�T_�0�l�|#i�ﵫȚ
�r�K���^�����+r�������e·.2�P���s�"L�>k��V:��0�6}Y{�n�����
`z�����f����lW�.��')c|U��&�BU%�y��S���Z��[E�M��ΓT#�9ay�{��6Ũ�.`��:����f��	��U�>7�j�\������X1�5͗@�_۾��_tn�s���n_\*�1{�� �sw
�.|IS����n�9�I:v,m-�iA����Y��anH��<��-�
~&9�	�:�@U;)�"/i��P�(tt!�����J�����!�a�Ս���$��ɪ34�h�~���NgC��>ϑ4o;r�{�Meb�ެb����/����*ڭn��ܖ��KWF:P٢|�{-��9\�n���C\�?��A��ڜ nBoa�$���J�~a��|�����͗5&ff�-AD{�Z��2hx�	Z�gx#���V;d�����WH�zڃ���ڒ]ђU���4m\�C��S��Ħϐճ#W%��% �L¯;���#�K=��&��/u��:-d�F�IY%εɾ��j^�(m�-��%�~�]p����,m��Y�ƍ����𵔲]yu絔8���(�m�dԐϥ�c�,6���;
ԙ�0_X/g�dqی���^@l��!���)�R7��Z(��N��j�$�i���Qh�9 ��Br���tɲ��ʖ��ϗ���ҌA5l��A�z1��p,����Nw��� 0��t�J:@u�w�o�8���e�]���;�-�޲i<�赗TM}��I�y+D��ׯ�9C*�n�=�ܰ�\�N���|���^o��Mc�����/�s>GNr���,(M��#�����;|��5h������R��3�(0Et�i������sNHF�$u��#ɫ*����1��bҚ� �q."��oi�:��S�r]#�], ��o_��7����wH�P��ա��h����9�pl�����a�������8C�5��;��UK��ZWC�%ަ�+�8�3�R���E`�8� n�Vw!ᆁs���#�v�̆�܄��>$G�H�fZzCҼ,p�����A��E4��攩*p�/�(]�W\��]#���<�2
z��|7(5&�{2A�`O��5&qdĦ�|]t>�|�ln�K��(�>@پ9��YR� I����[*-����!��$�S����W)%�4��+�sw�z�ڝW|��x]�^^�����Y6�K(.r��ot�D&d������.�w�^}68Dq���J۞�OX��N��Y �c-��ǻD�[��-�����p�Z���߹�k��aZ�����Ǔ�
�W�� p��)��ה.5@�wc�Q}	)?����9%�5��M��΅��"����7������i*YMwx�r0�%�`BaJZ�	I��I[��pY|� ʁe�t�}�^'i�ܻm���S���h�l�^ɘe�P^]=� ʠHQ�˓������?����ӌ��wB�����
C����ԕȈ�!�0�	$;�;�B���IY�~dE}�ع��P'+x������G����Ycp�M$j�����F���8����8V��z�cn/�3V˭Z�f|A��6����ƀ��S�0�9���Z�c)/Rw��k~��Ap�4ڑ�hI?�{�6�����V�®��[��YY�&Yv��Ph��IL�F�6��W�p���n�^��[Y�oZD�}s��xLk�<�<�`�����0�4. ��Unj�_3H� ���l�&/��R`l_�ht������_��e:��Ǿ���i/�F�FxO�eE�[s��|���g?�ǒf6J��n�Y-}��5[�Лf���g��S#@񃹶b⒕��Ɛ���T
���pZ�؃�3�7.x�A��f8}n ff��0�t�������+�*��Uyf�[�D�,6r�i����9�/��߭��wD�,��|[+0VK��Ѥ���]��O�G	=%�|�pkY}5�gӻG��gғ�83��"F�s9�=<܂7�,�qeE����4ۧg�8���Ҹ!z�Ox/]p���k�,��%n��t'�H�Uuy��'Tk�I;�*�1� ��HSehJ{V
�0�j���lس����8�<nLxx��N+��?�"�N~�*9��k��Bɶ��)
�bUEizYdwE��e?"Z�/"q�]B���`�V8R��������{刣�O���JC^���Ԛ`��9�`
�B0��!�=���vt���|v/��߶���R���Tm�3�<9祑=iz��!�@;�
�(:˪��>�<%���>�Y���-��������3d�����FKOi����`Ti*�2*��b��{v���v��0�+�zTێ�k�W�G� -F�^1M�4����R���^lT5�`���R�l���+�2SވM�<���p&�ct�i��w�)��VW�QQcH�S�ْ��$JL֠���f�ﬄu���Ά��t8b^k!�X�*9Q?��6ub0Y�+ M8�1��y�;K6ѱeD�}ڋ�R��!%��w*�t�qH���9�b�W�
߿�*�	҄>�$��G�i6F�CHn��S�����xW�� ���v3y_�#��d�hk��`����Ӛb?Mq�ps���²�t'�%�ǩ���#)��(al�<�r�LJ'���*�>	L�� �׌o�	_����-<�B�FҬ�&m+R��{}2����>��|�g��
ȏ���6L"�jMr��)^{���_t��F�xZ���@��C�B,�!�GH�����Z9$����k���:�Dk��xB��fYhwg>��$�Fg�J�<�2��ݛEI���߅'���$H?��V�b�
�?�1N(5p�!��*���D��?��U�evѭlm��)�LxEvJ�jH�`#��P����7\���ef��1?��.���>B�x��'mEbn�� �?ҫ�$s��nEӓv]��s�MSc�?�My��;��л��ߞIɸڻP�:��bH�T�f�㬕h�R��I��r�Ʒ埚L����!�@�� Sc�3څ�������\交	X�o����pAW@��G�-���.E�wGbp93��Z!��ԑw��D9�U��cHot�G\^E����mo�X+f�k�
�.����q§�$w?"W�����P���/��Osh�s�}]���m�isX[:�q8AX��)`@�W��Q[m��/����W�.�v���ez���Lf�ӕR�"�%lM�В�6�92��k�
.ރK�H�s�$���V�z#�&����5�4�GR(�0�X����_���h����׌��#_�Z��y��u�y�Sg�"��컜,�gHҞ�tM��8��i�v&�dpy%M��,h����E7%�n�W�bd�V@�p��
����q ;;@cu�IOrQ<I��1��P��x$��I(�:{D���q��F�7?D$�0��6Mr{n