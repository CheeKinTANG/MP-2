XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1>�!IV�m)]���s�mR��R�!,�3��/��W����7M� �v��&�ȶ�E��nSO����+	�.�ic'm9����DJ���������ϕ49�[|)#�wJ<���I��@=�۸ݲ��
ڹ��ڐF9�{p�8cH�omk�P���� ������Y�Glu#��ͱ�x�T�=��\�;�1���m)[��``�#)��ހ���ԥZw5��9��gV�#���\���	�GCU�� ]�P�-ϥ���c��]�����މ$�-Ӷ����+u/zj�ᚑ�;�㛵�o�G�Bjnq���Wg۳.M��*Cp��
R�cd���`5R�sa�D L��t����r���;)��.�vv]����P@,�Rk��q��V�]����(��ٞ�=���rjͧ�ֻ?&l��B'�B� 9z�Q6�g��]z�s�5 o.1��f�$�t�b��p���A����O8)HIe���VJ���|L�'~J ���am.2���4�^��ݧ�/�x�cc�D�[	�~�f����N#��^D�D����N >$BA'�g�?��ad�B�S��-���
��;����E�3NC�G�5F=�5��h�� ��p�[+�:�>�Ug��oD,ύ������W/v�(��}��]�K\h��1�Ɣ�D�)S	A�Hz���-f�ӌ� h��c�pMc�T���wsL�e�\���s�vS	�5�Jmd��9��k�Z��%n�-�1p�a��������]SR�XlxVHYEB    3fdc    1160��{,���CT#ߧ��k�Q&�@��e_AoFi*�&�eL}��a��Z��kE.{�%�����:9���<5/�k����KF3�J��9���2��/������Bs�y�"X߻���Y��ϩ�,�gvS�:#?���ͥ�Xy�!�k6[��^��n��N̑�g`�~ʩ*O�?A�o������盅y��	A���^��Ҕ��c�*�_
��A�ܘ6�/5+�g��eR�����-��X������#|��@�f>qEnb��pz��T:c�HFN��x���\�ld�mU���/�CR#6�˄�V�;�6U%��um�b#\�,�iJ���g�p���)��h�ɔ��� � p���~����sP"'�#:���Vq�d�r����~t�d#��^�J�sw��4]xը��MM=-K�,=�T6·���- �hH?�uu�<����Z��Lh��ʰv�O�����Kn��U��q�|]a�o'���o�E �oN�4��Y!�9��H�3�a�Ĭ�6gO���V`����=�S^(�II
^hm%n���0Z?Пerq��Z�����d��y��V��;E{���?3�χ�R�)1)�����L�?������P�am�S�.y���l�FU5�Jv7�!��&R���=��3&�]�d~���5�׷�*�E�&�o�wNf�O�} 6)� L��!>�~<�1vB>�$+��F9���=`Ǔ���<%Šh�.0�˫�#ĎW��|p�jִ���~q(��O��o�����Ã���?��N8�x���+ZΖ�T΂RŦ
V����H*T1-���iЙ�L�$_�N���\���� r�~M#��}�AA����*�Q�x���q�-��<#}�<}�+C���V�o:4Ub��3�>qm;1y��xT���0½��<��E�
��1����瞘i�G�����jJ���ބ�K�M]ʂ":] �^ ��q���E���
�����o�����]�`�� �V�5I��V6�aL����%D-�:�[y���T�]=�A���F���δ
m�<���@�k��;\،Q�s%�hQA6��r�Ͻ�핚�ɘ��9|ٴ���a@��u$FIu9Ƃ��٨�)��w��̼�c���V��������-�\H�E��o�+eo���3�'iU}圷fu�	�ç~ڲ�fF���Ȅ��a���_�i|�]��A�G�~Y�+B���2]Pi����ʨ���	4�n>���L]j��K{�RL���s�����0]!�,y�T�
�H�W*�GTP��,�S=[�v������.G�nyH/(�^��{kn2���U���㖄K�kM��p���u��J�H��e�<��z���l�4�B�E�~�z�U6���}�f۳��K�v��i���o27:Y�z�l�>��;�W�Qr�M�SC	��V��WkO�K˖�,=$r���c�U �Q�<@hT<���T��kU�مF�^�P�\;�=�a�fG~�� ��[q���S��>�ur�~A"-�բR=S.~�g��щ��i��_�~���ļF0v*�E���C����""�H��e����8|X�2�p��J#�>9<���uk����2��R,MzCz���	�Ϧ?!K�������H_s�5%A3��ux�u~GL ����]�w���T�_�ā�E��?�I�k�����Sl������ϸ�����"�z/6�w�{!��{An�+��<u��h��xݨ�5O�F��$b�Ġ 'G8v�n���R�wxmH��W
1:����Q8�t�'���b[ƹ3$w%��o���L#��j��M�DR0yR�5ł̈����5(d��9�`O��,(� u����;�N���m��3}d�w=�INy���-΃�N����Z��I
��.Y	mJ{~���������K�d�<G3�H
���(��m^x�^�@���a�H׺sfJ*i�vi�1)�G8>�sY���Ӹ�+�&,����{��q�N�#�w��bϫ[��͕X��� m�ݳ�K�J2]��K��"��dU���F>k_R��d?5�1�8ؼN������~n���$�NG��~	M��ꅣ�u����E@-_�4�����Yk�:��'�W�Aμ~��ou�K�b�E��HG������4Z��Bi�FB�5��ȓB)v�\�@s�zA��a/�fUIY]�=�D��'���}'�%g��J>#hp��dS�.���r�*K�����CΚ�°���#�xZ��Y��kJĒ�w���zlx+�#�;�`�=�<��Ȕӑ��ȓ��! $T��~�e�k��h\��#�m�&������T�?M�2�K٦��/Y�??��(8� 7M���?e�Le��8�b聑��{|U4?g� *f����D�Ko�9b����Uk�VpJ���P���BU��
�}B�� O2v����7
����C��܍w�v�IoO՜
lyT��]����.رѯ�aOR����Յ�����4��� g��~��Q?3�"�L
~!�����Z�0�x˛�]�-�0Q�v/v&�{nc�/�ae~r�.9�9a�'�A�JT1�`r�B;u� ܷΕZ(��<��O��JJ/l�c�J�ːG� Z|�22���x���ץ�zL�)�s�K�����X
�m~��V��BǙ9�����_�&h��>���HfM�S~Z��{�E��Y{)�����<]_EL��(��p���&U_q	p�#�����F4��<4�"ù /�R��C��&�5��K����fI��F�4�Oǉ]>���܍e]�ը���%22��闼�!xC)�]�����5:_[�]Z{������R�������4�)�w�r	i�G`�ݢ�׽޾�wvw�L���/�4��s�3��F��6��1�w�6I�81�zJ{��5P��,�Oj��{����liF�	L�rH�Ek9I��n�����&Y�����$�eP'�V�Ȧ9��샅�6]7�<��2G�n�掔wL���� �qe���ç'Z��X!0a	����sb�33fv�g�c�^��"&Q���9s�=��K��
���V
��6�:�^M�^n�9�d�	,�o|��#�'����Y��>��(��-��*�&�"v���]t���V��Z�ZU	فC{vS��R4�4���c%�G4�,�hB:=S�\�!���W��չ��5�R��3��X�Bh�GN+lkb|�[��t�t0A,||�5�|C�I���ՙQ�y�؛�56柚�z6�wwt[�0��}�����"wM�����>��Ӫ@�-9�}�Ax�A���æ��H,�M�#��g����w���"�����|�V���M�������\�Q�Ie����r)���4�3J���i2)J��^C�"�����l��i8K��3m���}��^�{��==�SĐNNq}H����"�YI����qy�YE2��X /�
j���C 2�Ȗ�F�V�d���w:�t�&�����As�6�����\.����5��Őri) 3���ְ��MPw�#W��0�yg����B�^�pzd."uz"%�jV��up)S�+aT����~P�������q�>����~>���6y$��!�^�tn$�e�jǨ	��Ȉ>(C�Q�M�ν�߯�`ݽ��=�������(�|(f+�8Z�����0�5�n�F�w$P=�'����7ƽҭ�c`w=�Z���@0�UyE�Ѱ��k�63��_���[@ݎcom&0q�VBD����������fN��i�Xr�o	����H�Ws��If�9*������p(�(08�$��ґ �����ce����/d��l�������.H������`���;F ��x���ͅ�Ie�J��.����Ttx˫�87��V̛T���P]ȶr��
ڤ'�����i�@��XF��t� ����L�[������*�}{�����;���
�]fJ;�>�A'����P�+G�7.��#]�qw�	��%l'�Hy77M-E��V'�ן�	D�^����.'U	�3M�R��r�\,r@V�F�0a��`�\��>�?�%��_�xŝ{�F��]�c|�BDX���N��� �t��B&��M):i�%�Hʒ��{zb�o�IX����W2Mq��rϱ^R��F=��fy���Ҩ�x�yS8��R��,���x���-=EzY�c/Ť)eƋ�z�pϘ�Г-��b���S�%��y��uzP\3
�δ5S!P�:X�oTo�'�n����:;����{H�{~� 9&�߆���t�00u�U����S������W����kC~|���.dWQ�c����^�/�;�'Xc<�,