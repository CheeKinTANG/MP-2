XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����KB�A���{��MJ뮖��6�a�BƤ�Uo�:��Il�_�*L$Wp�_蟚[1���B����7��	�=���*kt�����S��і[^�P������.����E<o؟+�}�L�r��U(Vߣf�W��&�1��$�9̋O���KuZnP��9I��G�dG�u�`�{ھ���3+IP��	� [����^B�D����P2:��`f�c�1[ҜD�7�
��r����� ��� 1/����I{qu������i�=ߖ�~��.%]m`=1�_���X��ʢ�Q������cK�5�q��Y�/�������7��� �O��%�_7�U������3�?�����d|j#R֟�G���+�6����\Tj��?;
�Z�ǞI�oo7S�A�!�k��ɒ�w��˛�] Rn*����I�u���hD/��yt�ڏ��E�1��߸g�<����4�SK��S���6�w�Wlp����kʸ����+����q�^:g��rׂ�2����\�ȱQ9;<6�v��@�}���QLL�~����%C&Kd[��<�.� ũA-@D9��`�����YE����[���D����߶�H�"n�h������qi�����@~�1~�Go�Lr�=L�B���~"�X��h���O��������hG�J����4׮��i.���|	8�U���n�v:�ͧϬ2FhvbC�
�T��H���#0�\�RPԸD�P��XlxVHYEB    3e93    10b0�t���B+��[�z �_�$�A!B�c³������^@E�O��C&��`)������c:���$r����
x�&6�D���(_��� ���`h�, 5�S)���i��,%�G�����Q2��A�]fz����c2��1�º1�ڿ)�q�S�+�1T�@�Y�w��^��_N����P�`M3�l��Ӥ
�Uf7(�w�|�˩IU���Mb�L�3D�o���� -j�qY��kP㽸y�
fTb����g�i�\��Wա9�t�>5z5h� ��0��@�� �C�� ���
K,�S���O�OV`�`�6j_cg�9�K��ƶKGls�^��J8����dK�ހ�^l�XB����>4��لD���8g�Z,&����PB��'X���f��K�� 1_��	4�ڈh|� [)�$�Ǥ�Ea���F�3o���YչJC�v#}�l�'�倇i��9�]���C��Z���G���Y*�sFp:|A1'+�o�����'�}
ƭ�YV�I���''�5Q�.�)��k�W�nM"�p�?�k�������& ��%C�h�5,�V>��Wc�!�?	����1�}R��a׷�Ǆ�EdS��{`��r�l���Z��a�.G�*�h�\��|.�8������hL�Aƻ��it��J�������h��L�HB��rb�#l"��Nw�
Z��g�Ho��,�\�ey��J�RQ���D#�xl����N�eoP>��ĉ��u:�8�o:�Ro��FA�ν6����Yy�bp;���j��0��V�_ 5rFيc���lg�^�D���bϰf3�XTd��W�M�\���|0��i�nҁ����:Z��W��up�z,= 1�%E����Q�}���"�[:�m��xÓ	د�da(+��G���a��1;Qqz [.9:닚2�,�3)�"��U>@Z�.�5&�id[���0jx��h�	Pr	:�>������_ۂ2R�H.�JW�Vā����S޷�CA��\�T�� �$[�e�# ��bs��f� �;��/�oH��C��E{�Āk*8�LgM�1�2�ܳ�W����X���.���7�t>1pg�ӿ8瞜ʗ`v���4zR�����Jle�K�*-���i���q�:��ڡA߶s0�<5h�BkAy��(�<��<�6s��wc�\JX~O<�|Y�{�
 �9to0N�*�ɰL|��B?y��k�b���KA�\��A�{&�b���쫪N` '1��_�IN�H����Ͻ@o���Z�nq�� 3�!4֣��;�=��@m[��"�DZNoo~2��ʎ1Ae�kiX����e��w��k
�:	�uk��5N6��HV�TR'o��^"h�[�a��|�� աS�2�V0�Dg��t����Z�����z�#�X��0I
��G��]���ۧ��5J��KG6/N�&g������ꮹEq1~V|�.2U=������dA2_��03��ʐ��3V;�FV�(%QG� e���[vP��Z^��G5��\�[���Y����������k߻Cz@��/hG�k���0\T�7П��1��(D��U�den�W�+��{�y6���.��a�D~��:f��M4��?��`Guu�<=�I��mJ�`�iy�R��bX}"nJd����_���c[�l�m�vч��d��Yv���� Z'��nuɁc�F�Ɨ��[xa�`�B�k�x݁�1	���sb?����"J<�SBF>F*;_u��B�h�y�^��<��?ƹ�}���*F�0 ��^.$Wp�j��"RVԖ�\V"�|^�)+����q����w�:ќ�Z"�����,�Q��/�5<˱<��2�s�&��J��>�^Ɇj�'�,J'�(i!�� �fk	b�U~��PE���& �uD_���$_]}�8>��	<��k�z��D�?�����|��AOXH!w3V����>�_r��QlH9]Ƈk�'O�6��߽�'��/Zo��n!���lAVR�H���k��9���25�^/E���Gf����"��no)*y��(+�|�d)��k,��X�ҷz��m���|0�}	Վ������-�f4(sL��E��ĕ��E��[60�g; �ǟJ⑤�����ب��gwde�l���v��4�.Ze�<��g)R���CkUU���&.����KGyk@��mk�v�ϖBb/�X_�l�i��9�X@��Έ���6�v��������Ux�)T���SI �����Yf{���?hp*Y��8���ϓf�	�oտ�Ѹx#�/�
Պ��h>{��J�n���cG�0������p8�I)��Y�.��1��8�����6,˹q�_N{+�n�x[�r�e����>�ɏQ֫/�j��ڝe�ك�G��`��NA�xt����!���T?=��;�3퉘tU�� ��a�+�� �EY��\�����>~���2��4�'ӣU�6��.o_5�J��[���z�uq�Zk(����o3��h���[7~�\�Ý�-Ϙ��G��h�j���>�T|���I$c�&Lޜ�As~*����_����涟�E�B�dB�A&��U�#�>�8����eɑ��`�9�q��y~A���.�}tCr�pܮ�+��2���F) ���:����㵜��2\��h��@�$/o8*���K�H���*6QEH(z"��G���>� pP͌ߑ�q�6�5.�:����=b�l�k�6�'���I�LV�:��	�B>�*��YE�KW�����U�Ŗ`���3�jx��J�俣R�D�AH=>
��i��-���׾?�/�]���=\'�����5����b.�c��4=�x:�G����W�?u�Z�]`>h���8t>S4��b;�x}Iq)v��ܢ���˩ofvA�a�A"�W,_�ͷ����j7W������)E�pN�e���cx�)s�z���姉����1F��$�j�F�.D��u�Q`�h���K��T[ft��(�����C�����G��3Yx���03\+�SR�ie��8����2���;l�|O���+�<�?Q�q�7oD*���yi�o�j�>l;�ѿdQѤ6,w��=����{��8t������b��v�%���'h����4�6e(�w߀�`F����l�>i���t�X3uk�w7���QA	%�� �Q/-� 8������ɧ���apk'�P�<���x�L�S�Q��i�"�����&��)�9M��y��U��������G�<iRশsPn��PY�g.�])+������jٗ��,�b����3Ε�_�T?��>&��v��l��ٟ�$��������րMI��Wqht�6�W����@�r�?^'Ng��*vL^���l��`����w�o"xt�o8��B�|��	R&ea�V��V"�]�1�`��H啌I�(�9�o���U�!�CU=#�`�rƯ�#��?�۪tE�F�����;�lZ3�����)�sȉ���ҳ�T$,�E,�ÛZ�A`f	P�x?��z5�e�5̅����[ x�%��JnW=3��u�w�䰄��$Ɔ�L!W���z��2\�f�^��W���I�;ٳ���I�"߼ZZWP�ޒ���A�<`����諫��师ӷ���UxA�N���/9J�_�K}��ߊz��$��a2TT=�
c�X�%_WH����zG�r��\if*�w!�<g,����5��A�����5c�zd3_k׃��Ny�R̉5�x6Ae�-�p'��5��)�d��`"g��j���ݤG�^" �_�qN>>��aE!mg�/��r��y*H�=��cg�����(�+����>�Ppqq�>�x5�/���D($9z�=�#�E}{�,��֒�H�(���R�Ƃ`�����
�GU@�#˜l��J甃�<
%!w�M�/�r��qiN�����;�H�a/�� ؚ6�_�e�/g���X��o?�f	�v�R=a7��j��!գ ?�0���u�7kr7�ON�|�Q�B��t}"/D��Ll\6-�ڍWj�-3�iː�}x�E�U`Άj��KkʚuD��:r���`sJM��?"�Ȇ��f��>����X�I����y���:�+�0х�~�Ǆ�dI�ۄɬE]����ni~��S�>P��ǟ�w�-y�:ml�`��q����S:���=|K�~�1FB�m������@�
���E_�fT��}�r���