XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������Z���G�ȮǄ�mm��PRV�U�V����m
=������Gv���"4�+���W��<������` �s2�n[o������8g��w��,��«_pmrC��"
#d���Z�9�y��O��nHr@��ߟy�Z���I��_rHñ-�oŏ��M��4� �V�	���R����ȫɛ$�~���M�#V��k"�s�@��43M)����<B��*I���8l1����0�#�Li�-�>�Y��6~����C_�p��5J�,Gf�*q��d�tPZ�UU��T�?�L�+���=<2c�[(�9����CoP$&-pq�Sd:Ӎ
o�h.-��k�|���^���y����r۽
d1��r2��C���q��B��5��ٯ�֞U`������Oy3Y�`�)���������T�+=89��7a��U:�.`�6%�)��v�lh���z=	}����:��P�MrA��Ip!X�x^4�va���M����"'����nn��1N��OTBl���ZCe�ޖ޲y\b���pWQ��4����>�z�}#�����w)z����*����*��f�-��ӇCӯ4�yHM��Zk#Qg�]�5�$�fQ����m�Hh×�gI�15F�4��hg��J�j.����&k��zM{Z&�T��"CH�	�_0%��o�o>�� �l3���+�ƪ���hs�A�<iU%������ ����:H�x>�I/�$B+OM�.3+E���%'�y��N�XlxVHYEB    fa00    2040�����/�_W��t��*�1h����hיf`��/tL���OW�mw	W�#��@�Y���@�u���AD���U�8�y]~����%�F[�0������/�n��e��m6��c��ȟ\Ծ#�X��e�΅S���x/����]ȼ^�O��5�W�?��x�1Qq6*�z�<1#p(1:���E�-�� ]4�����`�&T����5��e�����k9O����]�3�|\<������qF��6��>_S�w =x����2?�u�zz���Q#�Z:��6�����P@l9vK8�� =,���^��^I��w����%P4},S���w����e�,�a��l��8�$�����⋬H��͵d]����Y�����h���ص�����q`ae���78�G:���(G7��K�	I�d�9F���A��%ӕY�m����9��'�%�yi��Gv�_@��'u�J鑮��!:	��V芌����ړ�!���m%��$��a��������v��ʹ���Q�uiF�Q��A�I�S׷	�Ƽ�3��$�N-/L�õ��VG���%,1I��Z5����t]��yc�/3d.�Fm����~��<���:�B#5'[��[�zA㘑��0�I��ʲ��A�>BᎣ�$d��<��t��H��L�7�w�=US�#�p��Cg��F�GX*AK�[���:���I@���Vm�'WS��zz��D�'������=RC�V�P�G��-(��\^\�z2�8�E�no�7s4����n}��Pxu��u%v�n���0�NGtD�Ə��Jf�׉�[w����O����4���^ �Y��%j�
B5�L�-^�h���_d��jjGy��%X�L7�����[$��a97���~�����B�~eZ\'�XS��	�G14���(���*ľ��CИ�ǾxL+Q�XKwP[6����:���#48��KV�[+;6F��w�R?��(\��ȗu�Yk�
�k1b�0 �V��,�Ƃ���������h�!�܌<��y t�A�ȝ)��y }�K�ċ@4��J
�fT�^��	p��(��-�^|H,J�p��;�u]�d%�2�{�cSu�L:�)3L����0�Y,����p�����Vo�h��c��:ؼ1#�̈V%�eW{���zw��+��L& �GGɿƃ&̚K��5��9 ,�u��u?ɒ>`*�'�8ע���)��^9��P'lW��T������yy�U ��s\���1k�>��C)C����.�-�v@p���3�L�a�E��\7���ޔ�͈΋j���˸����
���ƛ�ۛ)ܪ��:"<) z�C�"��B\z�,���1� YpH��͎X��h��p��˹h6��
w���JT����Y�[l�l��JI}��̫G���W�|�TI>�Y�?�g F��������	{J�O�I��(CVy�W��p�q>�Z{݄V��1�*�v-O ���oLbelJ��u27cc��D�����<��Z*�R`A�hs�pO;�|�<X��(cjK�6erB�o*Iҋ0���ĝ,T,h)����S �6�:���G�'
�.Fk��{��l�H27c�~EXim��pJ��C�|��u|����;���*"����M]����$S�BU�Î�&�ie,�Ĭc8�������Ee�j��X��mxV ��#غ��6��G)��LZ�$ZX��~ �=�	'�h o�o�{0���6D%SvR�M�U��K��Ɓ!���\��H ��'!F)
ⰶ&��!+���$�?��ty��~����������6P��GQ֑����Y���6���8���R�Y��f�rFV4�r���]hо�30�Qw>Fw�0� L,OB/ހ=��(˯�9v���-��V��	 �޺{H��L�+��k���).qhWP�޵M(��z^֪E�T	J=	���.�F�=�Қ��6c�js�+�يٿD+�+���꤂Ŭ9�9���l�v��ɲY��\_-5�P%c��]���- #g���>7��	<����:��a��#-�7!�e�V/Ȓ8?����f�����
eX	w1D��"�0�̠��C�2�����^�.�"fϲ=t��
�p`a�8����V�u(���<���U���N���8�i����"�կ9�����p���t܃�Tg�&N �P�jb������DO>�a���D/\v���9�g+�:��.�$ڼ9ǳ@���*�R�ْP�w���H4�Oq��o��"w'�	���,���#.\-$��\n"��FM	��ˇ���m����vI��f��1:��S�An�aZ���K-RڟT��ub^Y�[*Q;�p]��Wl��Mc�_��ry�r�9�!b6f+3,�#�
�և;|���ᵴ���;V�ɢp���;Y�Kg ��KR�Č�S���[o����ȫ��az@-��TPd��3J��%�uY�>k=���Ր�A�� #�X;r.�k��U�q�̼ Y4�nH�m�A�'>y
&�����
tj��+<4�sK�q����R.}Q�۞�)���ސ����a�\�Gh��F��k,��֠�U���mG�n��nd+cX�M�)�^G��^�c8����@m��IaKܓ��L��ѮR�;�
�.*uh�(��ӯ}9ǲr\�#�P�T0�}��1�#�`ұ��S��!5�]2{+���p|���N,C���GF����w��
��}8�+̇���X��Ua�CFm���J���P$I���F���!�T����*�S��E��i�m�㙬M���v�@r�U���c��,�?$�İ)�V6N^�Ԟ �k��2��A��M\E5F�ܖn�P�S�����g����(�K��)�ʒ�GɊ4KX�<���l��Y����&U�:����v���^G~�Q�Q��3;�=_)�Vm���$>C%d_$�7�{[60 B8;�M
��/|B�L���u ���Io-Cߑ�2���rR �=r���a/(���_��x�d7E_O�!��v(����4E�
B�FQ�c����S��Ԛ3��w�E�ل�1}��<��r�Mͧ+��)?�� �����f�\��ʚ�n7hπQ�i����2��9 �HVH�r{��4	3��'�9|�4n���^��nO|����	���_S�7	1�Og�i�ót�8���0��|�i��{����Cwd6���}�Q�防�C�귀I�N=���������2^�P&{: l�'X4"qt�?ЧEV���-��f-�����a"�����^>���d6�֠�IFm�0��q;�����J�C�y�ϵrWf��l����e�pȘ�W>ig��a��4D��t{��3��O)�?�??!0'�ZI�UN>	{G*�򳪕W��=��H�t�v�e��9�\���6&��dp�l����^\B!́"Z�o���xM����ܔ(��kh@dq��?Zk����!ai`0ۄ����Q~o��h���F}O��2^q)Ei!-όE�%%�������f���sJ�(�U���F�B\H0�ȫR�AX� \Z��D}O�c�3�I!�֝Ԡ��h@�ҳ���c$2ZX�Z1�t��0�y�0�n�É?�!�lIO��.k��Se�QaRP�H���;��&Jo�s�>03�:��g����*��+�tz���<#�@MMe"ߦ�ՙ"a��.�i�ޠ��<;�s�+�MɖZ�'K�P��1��\I�e�Y������!���ˌ�ne.��13ħ��u����� e���x�߲A�JӋ)�{ylty��]S������� V$�����h���G��w#������Zu��*�R(�e^�/� T�hr�'��$�:'�����!�w^ �Z�� wp�F�F�I7�Z��{<3��6񰜓M#��s*�c�5 D_�x1�3��I�* !���RJ�a�C��O�a��M}?,ܑ�x�:�;�vd�]bB��<�r:�w�Mf��631��`���<I��m-E_Ձ~ϲ��;���^��S��1�d�$3W��Lݎ�#,0Q^��r����k/%*E��_9�Ez�����E*���"�ߠ;M��ni#���rW%Fp���T㍋����|!iB89O��'��D%��"��J�zQT��Q?�8D��9�𛏚�>�U�CM�̾]t�=P���m�����Ɩ���\��0s�T�7X��xS��Cݮ�SB�VȾ���v�0�:�����i)l (lq�/�?�s�:r�� ����,�fY]8�0���KC�Q�F� ����S�j����~�_��%s�;�vy��I�Rjw��`�i����DVz�R�M�~&�������C���j͇�����,�B�
t�k�f�f���D<'��c���6=z��fh���0���"W�*_[�ʵ`�V�V��+!����L���)"�G<>��(7g �c���ʠ�B_E�4�	�;�SR!LP��r
�Q}�I�&>͂����'}͐��}>���~��� sܿJ�)�}I<̟4��c�Y�D5�g2�&
�O�T,'�H�=u�ݕ�r;����}q�G��Z��Ӹw��̺�:����:n��:�Ț�=y_� ��1s�j�m�+��4*�����1s 	���:v��D��/���@t6qq�ROّ�z���aC����_6�w���w�����A"��V݀_M��c���N[A�5����<�h�"���s�o�=�	�ǭ��-�=dڒݚ��p'd�=�`�ПO�H�
'�����C8K3��*F�Zk)6�3�*!O�BG���A��vmč��m�=������r=��ފ�y��).�X0է��ɽZh�qU�UR-A��$�N�E��&��48��B'T���D�<��2H��l��>�Q���4O�_�K
aӱ�I,�	���p#���"�_�DuS*؈b����N�F��6�B�?_��J8xЙ2NIғ����,v`g:�Z��V��_�7j�-b^�$�d�m�!�@?(�=���%Ȩ�04i�,#?�Iu�p�n�[�ʄ2.0Mڶ��;��4ʴwW��`��zӨh��,A�)��Â$w��LM|�فn���Gƹ����[�	�9�/rUPJ*���x�	����"�Lhĵ�����H>bO����/�r_Սg�3�c�Bd���&T�X"X���Vf�����%�ڤ��r.��cU�?X�Z����{��#s�Yc��_y2��ȋ�]e^h��JW�y�j~��a�;�"B����M7�˕N���m���j��_�U�"N�)��tz!h{��c ���m_
��;�ט������xY�t�f8�xxU���d�3�3��=�K�*��y�&5'�/n�n�d�F�i�ؤ*��)��DNԗ[��;�Q�|���?�yr���4>���`9'��	c�L�!*o�8�tB?�3/O�C�q�d�C����J3Gmin�uw����!�0�g����#zD�I�7A������HTB؅f��wHˆ�<�o�2#@Ǚ���,��a�~wv
�%�����&���!���se�b�us�TW�;���~�s�a2}7�3u��Z���դ'����=�"����k`�˪�;�c��X%���=~5D�6ml���ﺹ���PO���x��9GG��JG��W��pR�p\:������}�wE�����%9:N�(�yy0jJ��q� z����$�q�{uD��68T���g�����{7���Os�!�̧�� �3�Q�v��w��MZ^��JL�^��Tv���`�ζ��O�e��L�1L�U�`����w:d�}��C}�g��y�˷��<�c ��)o@8�����#��u�*��66�� ��M@[�\�����DS~�+'��-��<�����<�Ɂ�	*Σ��J�B$Z�v�ǲ&K���T���L�G���!�<��}�X�s��p_8@�źI�${��׵ Ȕ��ILr:�R�̎Ec����i�����2έ�f�9'�@$��{�(��aK`���C���kx��ԭ����'ꕳ����r�W�����FEj�q�dT0��:��|��
��!���
1���`%��
p0���T3�7�.mu�u��؄��D��6r�� i�|��ј�SP�*]�x������
�w�?ɯ�����֓���H|������=tp	�I�UF�^�[:x�q��@�h%y�*R����S����IK#�a176G����w�B�-̈F�Z��e.ģ�V��#�U ��% �����r)Ȉ��x�S9����`?!�>��d`�o0s�QwU�1D�~�3��2I�.pM�aCw��*�b�d�S��� �;��ڿ�������y���[~�h̰Y�PBk���UU��.l���R.�%"F$�l�9kvl���Qf���I0��=۫@M�1��M_ � a�6��4��&Bb��-c2��8gsfzt|��O0utv�Ic���B]��~[`Uv}��Og�DJ����{��ˀ����@��sRr�B$��3?c����}7��$ ݙ¨�w ��c
�UfWI�Kq�#qu��3�u֊������N��izdظF�37�4��W@1>��[�#�W�)T�f�6�ї�(/E�qݾ8������]�wȨ1�J7��w��\~�7�^m����o����Q�nG�e�sb�.�z���pd����M�A%-(X����k0�F5k��y����+���.�f�+̾�1NS��,HԮ�����V���v������8�6�H�И�x��o
�k����?��-���iB�Y&�;=��l�؆0S>�ZL��5ıVK�:/���L'�b�Y|J�cfY���L��U��(���?QR�iv˵���N�M�Ȑo������25Ӵ�P�s�h  3c�qꮅIn_�!�������>!|�j%V L�2GJ��2�5��P�b�&0J�q�ؕn�Jȝ®�{�*�n��G2��zQE�������o44��1�c�[�N��#�_�(T(��7�J����uF�U���Y��@����L6�|���u@�Wo\-��K֪"�$qڅr�Q���x~#�������y!s��9���`�&?�zO�M`ӟ���;���U�c
������ �V�S��Q��_��rZ���I>�^+���] g�6:���;G���G�|\�^/��Uݸ��6*�x�J��_��	%=����
��t�~�ĭ�Wy�M�>ƶ�$ŝ�<��_��@�mJ�;�Ф�l�^P����4UĲ2A=�'\${L\��I��&�_;q㐏=o��� ���u�(q�Q����y�|OMI�e|�`��u�9nJ����>�;�W[���4�?b�� ���]�U����FEJ�����g��
!�i�����/��J|t��N�0���tǈ��p�_��C���|n�
���V�x�w�6��j��0��Xe��>��S�X�m]�oYS�)y%P\ ^D��Ec}�p��!�j��l{�).��xc��ql7��8n���+�O�slw�34��h��\��ׅRɣd���A�ͬ���N�U/�
��<RU�i��_�45vT=7�1m��K�G:ł�%f�p�X���;��u�=��;,U�b!C��Pu�]7ON��Z�7j�sĨ����d�K���o A�he�(N���_$+"R?]1������	�������{���TT.`��M���R�L�1�u�ګ"��:8U����ER^"�Tcm�l�ޯhx����˱�s�_� w>R���4���1e'��qD�y6Aw�_jH^��h������a�u�x�.�?�����J`Q��V�I[��_·�<
��u���AT!���XK�X����g���`��ŋ���+��,Z��dsӖx��2{l&N�~2,����
��358T^̣�9�&4K��� '.gޝ��|W�V�f���ēx�?Y �i"���~�E��R����'��OP�Ɣ��I�b'=�Ã��ȝ�PD�gƙ:׈��pȺ�I����}�x������]NnQ��7$���\`Sc;Qy�rY"~⇃���	�=6�Z5h����k�����q$���e�����u�[~�8�λZ�|���Ҍ���bfHt�tQ�5��D�b�V\1/���Iv����9�\��°H��%�I�w"M:jXlxVHYEB    4f62     b50ֱ-���J��@���[�U�E:�>7nR�ۚ�]rI�3$������)�����U0P��2�U�w:x{�8�E?4oմnݘ�$t�*)��:��ic��6�k�/!���t�v�`c <"^�� �	N�-�-�)E��^_��;Hт�.�\�Kȕ��q��h�]&��oS��^���: ��O_֔��U'�̘W���F��Y��2݄R�6�`qR�9��]�,�]�Ago$��1 �!zuQ���բv�85�0�k�/�Ҕ_�x\���4-�w�P,�m�����*6P�a+�/e� �v�<Y<ڷ<��W��ĳ��!��������A�f�ŝ�
%��&����i��J2_��DA�#�j�6�m�!]i
-����[�\B4c"� �.;~ה4��f����������\�I�P{ժ�ɸ����s�R-�y-��a;�u�<����4"=�0T�7Ffm]YMOԋo֘U"2�[>Ɉ��!�"�����2�?+�V+���GU#w�{룑8$xd�H�!���y�GF�cK�2.�P�̭MT����d+9���6K�A�Ln�T1C=u�\l�RFt�^����i*m�7��|t����y��~t.�g�[�C���e�E���:���_xñ3�u:C�]�8�l��شj��\2��Ybd�3���d-LcA�p8��%S8z̙��y���٠B�HkW����b�1`X��{.��}Nk�t�����޹g֫�ŠVU�cL�=|��Y%�Pq����;B1��c�l���OU�0Δ�W��#� ��¬�,�sM*�GF�:�%��h>��W�	NN�)T�5�N�[{�z�������p�d=G��$�G�|�B����G��Y�5U�~	%��S0ͰbE�q�KPv�f8Ph"�;�*N���MW?c[[��p�&[T�MU��nT�	V�+��8}�k7��ß������\2c���͜��u�d��^���3]�s�Iڗ���Cg�Nx@�I��VK��p�ٛ~���$O-��	PU�<_����&#�c(��#��4�5~�tF��D��#��p3�������pJ+f֒�.�{?����s�!��3�\dg]w�B�L��R�#(Z���u�jc�3�.��L���d:Z��%�j��K����6����$�;o<�̑�Q�
��1j�`�@�-i�p!Q���}ZXk��p�ɬ�v�W.�������o5�ݑT	n�P�g�
��w�Mߩ�0 P�~��q�e��vڱ7f�T�T�'���<p���~��M�����;m������t�B���cX\�=��gW��'�R6�4E�m����2��}^��E�n"��V�Rq�S$v��d�0��a��^�ʽ�K.*����\��`�<��/5�'(Af�KJxb��Zc��mR��
�T�#�c��Hɬpb���?A�#;�U]��Դ+��yR�X8��.��#��όO����ks�;�1���`�������%�%���R��E���h�����j�����&�)�F�^�F�δ^Y
/�Wj���;�R��}�~�+��eEuG�1B��[.R/�;!dNx����ZzL䉯�
G�D��|X����Y�����F�ڪ���� v�}_w񋛽oߏ7�-���1��{�gto<I�Ŭ����J���sٞ(��#�j�&m� ����D +���T��z{� ��|$�D�wbX��a$n�L�N7��+=@ᓰAw�n�}�0�ֺ���B�a�Z$���X�k,�{�S��Q�4�z�R��S+����aֆ1D,;��<��0z`��K'4o����\�Qd�][��*����aN
a�����N��2oO�u.�ƭ�$_w�5=j��kߙ��	Р(33DR�Vاe&�7��T?�ي�α���,�W\wP���PGCD~)�l������2��]E�\������Pss�����;��a �EF�W�9gT�o-�7����#�sY��}
����H�F��3��q�̏)6D'x*M�$�S�2MʉAjZl$^y �������өÁ��}�(%���H�xM<���YQ`�^ v��j���2.��Z�Y��L��nMf_��ɏ�w���������w݇�����Q�
O0��e�1�MQ�+�Ԓ
E�̤�OS:I��ծ���1�x��B���cZ�U8}^f
�k�D�:��g�O)\7%��YX�`2�iPwF!93�nv�m?�(GkTd�����e>:N;�5��W
sU�Z��0&�
m�;-�u<_�~�[�����dc���\]��ƿ-Έ/�&�x]|��ksY8:q����G�u��5�����5 2A��
�i�C㰳���USGm{�������~j9�"���n�mq���x@Dq6�w�Ϡ�����3A.i#Eҳ��C��{���u���Q��9;��%Qet;o��}��L����8�hy�
�k��*�9����7�?hc葝��#Y�R����|?���2��n<Ƞ�}��<�bX��>Sg���K��Q�+�:��j��>}k^�"������k�V#�Ն�֞��~��a	�^3�(�f��τj'+쌣�j�9_S�� 5� ��G��]~~�4ތ��B�Ï>�@|vJ=I�p�0���Pк��`j���
��F���=�ї�,��S��>~L��ֹ}��*�A+�P�3�%�>���K��:�#�٥�:�-�44�.'h)���gUFp�՚��6^�-��}�t�u��5�O���>��Yi��WtT
�@�&UT7�����s��� ޣ�p��ޕa������]��	���8 R�ϻ�DX��%���B���Ag�ɰ�>�����Ig���{�^�o�7_