XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5Ϭ[5���A�\�ҺK�|mj�V��1���iׄ���'ր70;�	$�X�S�-7�RIB���R�YR�E�?>]�EJ(̒�jJN����_[��QL��|Y��@ +�"h���¤�1�R�x�J8�"�B������m��	�Ϩ�C�����*=5��W[�]���w�8��;���&�v�h}�[a`<Q��TT�o�.B�1x����B&�Y��Ɯ��%�J"H*�s��r��ԗE�:0G���U�
��8���cG�ɻ	���d�|x��P���S�D��Yz-/�Y,�V�&�&|�id��R�sZJd��jd�ϗͩ8O]
�CZ�0:��P��At�tC��b����:5V��%_�c�����Y�z�S�;�F�1$��1c4�-h~Q���_��i�B�A���\������K|�=��;�kI�s�32�,��K�ڏ �r�ra����W�n�F�qZ�/�)?����	���ۼiRH�h{��[���	����{1$x�P���?��"���p�S���dmfL�ϒ2��=��]�j��(]:J̳/����q�7��|&8�Ið�f�Ee2ҧ�7^�(���BG?��N��%�Jk�$l�?�.SI���:�}�t�*��@�ǔ�y���إ�$�۳o�٠��#JЦ�V+V}$t��MIl��S������f�.�l��X�Y��͸B~{
��8���������i�D�B�5~��l깭H�#���r�7!XlxVHYEB    9fc7    1fd0.��J�)[=�o��gQBv�t�)�_*���c�O�:��N}!+a�iVW��P�6�T�N��\��Rd��<�/|g�ϱ�k�N'p�\�9=�\�Q��-|a4���'�Ca�ub�&��T�l�-�{�*����3�S^�\��� �S'K��*��f<�j����>����{�Y�=B����)Ԗ>��媐��1��UM\1�ҹ�x=���bo��'�*�ί4��I(̯f�Ƃ�%���c�v4���U�_L�h6������kS�s}�i*�T�2�z��<C@O��| ����N�|�߻`��dS�����Tʻmð��jn�ae�;@߀s�_�5N|tU���gy=|�lp�]��o ��֍*�r1VY�fZ�:ƈ�d���v�&$o\�!YҥR�UXS)+w���go�s$�$�[A��%�L�s���ʰ��,Rؾo>���5�]7�X���24J�Y���P�'͹	�h�=l�6}��oax;���g�>�~�<c	�@O��:�-?|��(���,����5х�}���}̝=�..�͘�.Z辺�6���ar��).�#���K��ĉ�-��w�:r��+Λ�{�d�5CBrdt]������&%F�f����n{��+�l��_����);�o?oh��#_2q����0��'�����pq�{\��*&-�I}�C��`��{"���*�7��O}JOesF����7 ]C��^g���) �����GZ��)�����V��2�>.į<ߜ{6[� ��e���o��.��k�[�X%Vk�9~^��v�+Y#E����"�l=�8��-R��<E�ǻ\��V�O�-�I=�yq��	ۧ��Pd@��=0�AO̼�"V��|�3 s>P:jL�ͻ����p����Q��*l�DrO��Q�[��)��2`�*t�-�+�1vI��q����fs�Y�b�Ɂ�vw��&r�y����`��Ը@;�&yiG��[���C�w�O.�����`G^pn1Zx�����[yK8rn�t-�"�������_��TXEh���h2��X<ZZ��+�h���n��B���P@�>�jiǅ[�c�/�����8�����Y�
�)��B���*N���\�%����d����Ktª� �Șq�u�^X�k�C����ѮY�(p�:&��9t�irz��Pv�T>�{�y:�-�� ���I�]�9�5D[_8�R���O����\�=�Ak7�}.�����w7�������<gK��b�/��ˤ8+���nD��J���[#�<w�e�R9���u��ؼ�� A�|wӸv�n�[�+VގЯ���CA��)����_����j�͎�FFE�4�>�g�-ml�&+���� ��h|�3����D�#z͊��n[�����|��ی�.�������4�&�FCވ��&QξnN����Am�����B���T.�Z8t�Jj� 3-+� ѷ�C� �J��m�Ӂ|�1g��?ZL_�9�zEK1�<O�oa�Lvϯ��YΠ�oԖ��H~�5�hЀ��Y�'�l�U���s��f�(���9v��^D#-������l�ǋ��+��� �lO��J2C2ԙy���d-؁�b��NA���� -�l��#����8��I{��?��V]�Qz&� �TƖKAU�8��04ξW��ՍkG��� ���=(S������Q�e)l]���}5w�̢~T�!�!̲�˦� w��K�b^J�+K�����	���?Q���9zU��Q)�ό�E]�H�Lƀ3[M�:0�.g8��]o8�r8O�&����\#�L:j�kH�������
&����~$ˀ2�}��<n4_Ef�C��e�}h?���]V�N�i5�4����	z��
�(]).x������H�������E�N�a/	��o&W�I���*$E/�=4mP"�HC�n�L��z�-\z��"e��M��X�Q��NQ����;�#��~�V�RQqҨ[/��1��>��d5�9\�~��W��A��))KNz��+ K�g�yb�]o�����K�����|J�U"��;y@���8��,�Nv���������=�^��ܓձ��\�J� ����z_���q����OV�1�<�J�?x^�i�WE� �8�d���f+��M�N}ڞu�쫍�p�R�*�Y=�4��/80d!G*x�D?�%zi�jB}���ۋ��m�v�}��?�M��S?� �
����ڈO��.ӆ�$׶��y���fޯ�����s�&i1W0�-�����Oj��jK��5�Τ~��}�h^Q:(iK�ueȴJ���)�o*��]�(dS�{=��#zsy2I��q�hn~���Dҵ�W.��O�"}Vԭ�;� a}��W���mQ�ԁ�n�zם�w� ���2��A�p�	y�
f����˙+���r�����.-A���i����*gI#\��`'*ʂ��B�����ύ�a��Zd�� 쫳����Y��7��uk^'7��(���4�&�C1���<�z|G�oHL�8��tl�w��-�:�ax��4]��|~-�;W��<0�{`Ox��g�V]x�,׃�'�h��FO��cP����eb1:�?�0�sTcc,�]Ǵ2������u�x���q�0�.��.^���b��O�z���A��7vyr�*���-x'?�N�������N/�@�|4���j�-I������Q��r�+e���9{���n�Y��yFR#0wb�����7t�E�`te� c�����'Ah�6E4pT�����w�(c\*`�=�j�&W|l�8�
�m1DX�ഺ�x�M����H��b��f�De���d�=��r6��r�ha�!��~@+*4>v1���j�=#[7�D�Y椴z}��zS�l̠`Y!,ц��vbÔ��<�Ep���S�6c�i�hȩ\��^x1�8WIh:ӥX"�ӭ�茶���z-=���z��Ñ����QϮ&���ؓ�c��P���J�tQ�L�~��۴�D����g�-��F���r���z���(�]-pB���	�gt�[�.Y.ڈ��0R���ԭ���V~��^9Ӥ�T�!��hhA�n�_��H���M}��+ ��"71$�ם��]���� 	Q+F̙�E�GТp��k��b��o�����{��IJ��m���8K���v�<�m ��upҁA�m���,���G�3cW ��iZ��+v4�`�F�=�Sǌ4�D �|�89}�VL�7�i_�<w�s�y%,�1����	�P���1h����&��z�n]�,�C� ��J��Li�.�ja��`�|�w`�7V]�h*:��/�c�y㮍%B݁}�1#Qztꩅ�l7}u�[����Yd���`�j�
�Һ{���\�w� F�Y����_��2��DZ6��yF
L���ƲeP��~Q��H+Jc�|L{!U�N#��xe��p�i�2(�1��p�~U������W9T��%�<us�m+i��H�{,%�5�S_aw��I���W��ҕoA�#�&ti��c��.+ċ�-�K��k�4�p&�}��5&��m�
���8�}�c�Ho��_A�&����ܰ,@�_���#UP+3�<W��'#k+�����G�\��e�JQt�rHf͞���P�J6�'O��n�E��s��˝��"ƥ
��-��3��OS[	TD�fwۭcZZ Oϓ�8��.K
����/�[{K�V_�f�'
X�5���R8�lhzrdyyZ�x����]K!J����b�'3t�y��4�3�p�~+�Yi?�uq��28ك5�>�r�\��tE��+�qƅӄ<���ңu�А����j>���L����q#vߑ�m���{�����R��U�p�&�!t"_d��3��?���S�O#����j�k�zT�bs�]�%�T�-��Z+N�q�z!Gܰ@ƺ��t�W求 ��(ʷ�#bb)�i�:2���l�)��!Dd@]e��JMb�x�YT����J����bS!pV�����Bu�SXI��b�¬�,�n����v�P�
�*�����.E4i�&u���q��d��ͷOM���!<������<U�)��b�I9�vO@O(?���<Oe|Ԭ���7\��nh�S+f��^z��(JV�N�@����u�Vr�\�eB������!`�@����It'�Pń`�\6	���JX�+AIH}4��[h4N�ۯ�c����>��\�W�shQ�M$E�tfq�M�Ą��g�^������X+��O`B���/�C�����C#�=��%���y�{���=�	Np��W	��7�>�4�|�gQ1h���gO`�h�%��u�D��ܪ�?�Nb�
� �v���W�O`郴����2�J�y��$jٙ<���d�eN#M2�_�:'|FKm�{h�Kpu�p���b���}��4qlg�ln���yW�v��]�B�r����T��]�ݠ1H�
�����LQ��ku<�NRW�-~1�QL���xn`*�de�O$�lpz8��<Q9��A3v�l��Z[#T���yx:M0�c\�ќa������y�5�)�/H������L��/����I�:{���+6JEª�%և��OdVޘ�J�e'���r�F�L��	
�de��q��"@O�a�|�N����H �����>�E�$0$:�9J�|�aZWԋ�I�EzGD�����s���D'�$]7'�ȉ�B^�������A��8#������\^BAw��hsv�k�gZ����fgN�_���B�S8�G�H`��*�ף��o/'�*�ބ�}��/-�و�ԣ��1m������8;ܽN�ђ��-|�4I���Y0�򬘚��╜��3�R�̆��@T��B���B/*�d���?�[�`�=zQ �����w�`>���yp;�6_�s��olM��)�iθ��L��a��l����;:��}���W�V���H,�J�>�C�����X�9��V$�t�܁ŏ��+J�N�D��R���Db��n�ф��N��S�/�yO�������i����t`�pM�O�=V�>3?�s��d[��?�}�3����4Q�*E̍[���*ږ�3��
�m׺�eP���"ᙻ�ěօ���\ �{��g��*� ����V[���/8)��t�&��ê<�:@��6�����a��И�)�p*���&��2�J���b�B&ă�eiX��Ú�4=i"f OJ��ߕU�$�#��_���1����&�?4j��S��>%��N*�v��m,�D �n���J�J����lI���&��/��USc���g��(��(cV��� V*�����8�:%�@J����'��Y��:�
8��/����
�!���<��dS�x� �Q+5����s����ÿ���a"W�4�T�|�5U<�{ EG��m��/`�G�i���e�`T�	�_t�c���m�4Ƹ���#
L��+U9&z��c��R-A!�p�&�L�h)e��f.�\�ms���Q&D�� ���&��Q��]�e�q����=� �[�ծ6�a5���u'��>��X��)s�L�a��Cp1y1;�_)�ͻrx^��>��͸4
!�q���J-f�|}��G��=�]B��2a/��K\��^�� C��!�?��[�ں�^ȱS��ũ�����isG�=8�ߊ8��ɽ[�:ҡ�0h�>��n4wXYǞM#��'���fN�ڃB4lƙ���g��&�������|��71�#j{6�UGx�
��j�B͕��aX2)��P�eܢ�I��)�;4��I��j�	9���@֓�|�fIaa�N�iy��]L�EW8R�����IW�A�v>�1T�M��&�{'�a�`I�nDH-Q���zz�.
[�p/�rD��zY�@��� ]�JG����Z>"���i�k��'����ض�#�
3��aW&�7��7�3v��#��.�qQ̟�@���ѽ���=�N��I�m/wJ�Ik['j�w�@��t��d�{�ǵ�j��j���6x�2�m�5cFC��ON��t*�nȾ��k���ͬ�/CD�v�D��\r���F���q�Co\ܦ!�'d�2A���2y������OO���Tu> ��{A�I@��L�~��hOi��?�����A��s���@
��zU�D,]�cԓr���"��Q9b��XW/������ֱ�b��M�
�����*�i��ދl�!/���r� U�Q�=���(��*��1�E�u����?|}�$�v�s�i!hz��y�u���_P�Y ��@h�<b�1�%��Ohul����-A��J��sMe�������z[��e{�4�G��O%/�f���v1)%��|_|��,��pޥ~�B�@D�1�)���	4���B;[	$d�p�ˢ�Z r�BwAA&�d;fv`���jT�ɝ/A�K<K�o�f|w2K�y9�������kh�K�af rG�r��LƇ')u-nO�AnC�"��; $(�=��jⷯ�N
�#�`���d�}Fg����*O����>�PƠ�U�m<�Qp"A�Yo�Z�����ج�,+^4��
�[Ʊ}���U��j�e��Z��I��������63�ƫ�����	+�~��Ct P�����1�.�'hFdPJf�8q
4oۃ���-��2L^�t��<~�WPF!I,���:iҍ;_}E�������,1^���T
����dzj%���Γ\Z�f
�Zfx������ ;�7�TG��z)%�ϊ�[k���fBtc��o�B����yN��H^�N�AYа�|�IZM��^Pl=�b��Y΂����e0���90<T������T�K#�������1�!��R�G��Oe�<��詠`�k27���{G+`���j�w�Τ׳���4O=�����vH�R�l�L
����-𭞇w� L'�r�RX�׮�8�M��$seͪx�>��%��aaxuN�Z�u[ۚˣT�X@,�r'$ID�}O�l�C\~�+�O.`���5c��\����
v���-Jp�$�]�	�ii���CBǺ�	��TP�K���"��er�Ή$�%bK�݆��/�\;�	M��̳|ϰ�ɽ���;Z��I���wg|��m鮐RCف^-�D�*_+zwy��!eܧa����
��m���.<���$�q%np�War��Y�����%����ǚ�?�Oz������a���wJŀ��� M�(�����6m����S�t���.�	�ĥ�w�c�F�ffÕ[���H�@�D��;J�7HE��[�zjwǕ>�� ��+��w �Dv���Iܕj����Ά�
/Z6���q�`�����X�b3�,�hO*�6#�y�$?m��㶻�ud����Y��~�Q'�Q�1]$�v�oy�b�j!�U}�/m�ՕS���ރ���g̅]z��z�)�Š�|ȹh�-��ʨe&��/qgK��Q_�C�(j�f��_�ƻ|C�m��^�'�ē��D���V؝u��� o@��5�&���d�EB�R�`��۴��\s� xe�|7�gz{���^�}K<Ċ���[�dd�
�dM�C3l�ʩ`6��QL
����<���9���4���o�R�>CJ�X��?g.�~c0�,���b���e�S?u��t�?[2Q�u-	g��?��5�����3��[m��I?S�k�1�ߍ%[�o'��mԤ���<1�o2K���-eĚ�X�c�K��>����Ty�蛛PN�taIE�* �Rq"�/S$i��},�h\��@����]��78�G�-8��J�a%�m�\���gk�?,�b�n�|��%^��v�䐘ǰ���o.{�aX/L9+���������k��ax�Jf��t}	�Dc��ҳ��(��F�^H�8R���)����H�;r(|3Ow�N��Ҁ$(��{p�՘h�ʏ�ơ}�f[��J���]�!aĘd��Sl1(��B�\���6yu%}�z���v��M�Ѷ@��>��'�燘'�G��,
�^����I�� � ŊR&\q�q�b