XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H2�QɎ��P
H���TM9�����'��\z���od��������T��Յ��r�f@��U�-��1���d��dL�)ÞV�!�!W�إ`��F�Yn�l]�@�X��ig;';[�z/N&%s r���>��fҤ�H��N��i	�;�Kt� �Z���=��U���K�Nܢ�L�r��r��_z���<��c�|�&�)��=�n��yRk�t�y����@����WJ\����E��<K;���.�u���:̅]�c���� ��Ѩ�W6�t����Ÿ����	8[�����;>�J�O��>gK����A��R�O�0���H�<�9qD�B���N��k?� ��2�V�~�tj��KBū�N�����Uڽ�� �H����E��b܂ś���|H��BA+�v@*!G��>F���r�'V\��(r/ &��(�k��b.�)/&v�M��_$3�l0��Y#�޺x.�H���j�b�M��0@dH;��������2�`�-��
)���=!w����hxA��tS�⣸Ȗ��
�3 Tx���%G�y�$�#�^ +�	|���ut[8�����U݀����%%+u.y�X�M�����,r��放���vi�V���T���$��xC��0W��ɦ�r5�Ål���W����}q��"a��]1怓9!^���F	m��})�%�������>u�'۷#	�i��.�b+v�g�e���x�d�����n[�N�����O	���XlxVHYEB    3b09     f80�}r��Qh�Q��,�rץ��s��/�X�B�g@~�{čq%���C�z�O�P/��i�w۷$����/�C�TZ�.�=S�z+�Rp�Ʋ�O�jQek����H4:Ċ��[�� ���q	{��j����p]����=c��uگ��(c#b�1l�$�h�����H�}�0 �n�>�콙]����D����b�\Pe8���������^��C�N.�����'�f|�RU���ߪ������r�B��H-��r>���d�U�e|��4]�#�a�o���=��&�;<������B�0u�{>�ټ F_�R;K?e���w�Ǚ�.�m�����U�ْlm)�v�[�� ���#Bx5	�5�&'���`�I]%Ĳ\R%��|�]l��O.���|��9�M6~�!��3�j��#4�_��e$�?���\[
CP�:�q�����<B���0g��)̡�Ϡ8A��7������h�:���A�bA��`4��}�H��$/a�V�������@s���n�4T�T٭l����k��;S1���^�il�01���ѩy��9�V��*��ʴ��8�Q���r%ޭ*aNI�1Z-�jpO��&" ��𺹻ٰqK�
V�������U^����r	c��ea���e��n�ĬRQjK���VQ4P�%9ZT���E�Yd�1�,Vƻ6o�L��eӔ�� �f�<S�Ά�	���:���nf=a�S� ͢��( W�ҡ^@W��H6\�3qٺ��������dAGJمĖ�wXv�K����C�T�+�D���\f�5�� �H���%%��i#TO������&V��i��KK.�JhnA
f'?
�n��	xQ~�5<��sۊaeS� U'f��w��9=��㫽�'��JB$�J7ѓ��P�1.�>ғEr�+�nXk��ym��b?��}5��j��2�uG��ɗ��n��
�j��� �9ҕ�Qa�v�t���ؤ*�G���h�d�V�m�W�SB6��������g��U�&l�rs	tj�����t��;_ CU錕����&Xd�Db�-?y0|���"�	�u%��I���t$�E'�
����v�
l�=.)}��T/��S&G۹�)#��q_��wWBf2�Aȅ�Λ:��P;�;��Ju����{�����"�"�M�����+P�����h,�d�1ih
o�k����d�X�K���jQ���+�F�Ь?�!u�!����SZ����ᙝ��3��C��ϟ�e���g;���a� �ۆ6�Um�^��f^��N݊�oQ�}�?9�~�8���W�+�%��i���m�'��h�����;�mW!�_����w�S�S΋������\am�q�{�@���N������o���5���L��n���N�|k̔PH�_�K[PЭh|>	z@�}�d[�1�L�Ki�YA�蘿 �R�o���6�)��d�(n�
����j�-�WvJ��H����	�8Ԣ���]aS�*S>6n��Lf9r���_<m�4��|3%L��HBS��m4�w=N7<�=֨��(M�1|\��|{�Ӭl��������i�_�IlB���|+^Z���RF�T���J�������wp�
B�7|���oU�RtkB _��eKY�������M���zNi�O<��J��B1�Z3E����;� �I���� �mޡ��A�52������0��K<��О�3!���ѼR ����cz���#д�Km5����B#rZ�,�⽞ͦ��	�V�ĕ�����	7M�d5�Q}�B����Mm��Dg���kW�~�S�h�G\76~����-��z��K;rW�������V�y��b�Mz�y�4��2� C�9���ᷞ�d�n(�sy.��@�TXv�(�e'��q�NA-ո���&��Ӄ�zP��H�ş�^�*6��@�	��I#�#�KbӋ+>�F��&~́2N~��a�]u5=���*������"�Hzc>-��|�)�^�6�z���=������4[��-:��Zyx?ZI��yu�v��+�0���/u������|��}k��O��E�-�.���]�Q�d6ͺ9���� "��!n���\g��OT�$y�r��0]�+@=lsU$�ɥ���ʲ% M���F%Z7֬��ft����X'1*0:���(%g怞�U=w��q8C-�Y>�S���0�"���ܲ0�0Ie�����3�E�u��%y��.�Z6:1e��[D3���\�7�v��,x�|���7t�r�ym��Q��\���N�CN�_��e�L���P�6G��Z�8&{�������ru��>�`�ì̗��@7���*�ƭ�y#2Y���`)��i2�������j�v�=pMԨ�a�a���Rq�%]��5I֑H*��lAX� n�r7�`#$�	�8i��/K���������qa�"�Ył�"d�Z�|���3�JO�v����6A=O^���bw�m!�rlS�����?l�z+b����:���ЀV[�
����;:�������"��C���ő����n���L���]��}%es�2Sվֈ|��O��c|��G�����j�St -�+�_�q[-M$x^��fQ'��w���.�g{��6Ekq���Q�����vM�J9���l��[���G���F�$�4M_;%}ˈ\���rqڹ�ǣ�����ړ-���3'��J#X�/4'�+*mh�S�PI��%Ο��I9�)�������|bB���ش�5a"Mׅ_�|7�6��`���
֚��yR�6�k�MA|[S��۸�5�Hm8�����hk���� �SN�Y1+*��7�Y����xe[�,��l���Q�'ғE�5����2����R���@D�W(�X�q��� �2xI�;-��-2���s��A�Ħ}$�.l���T�J������3��1ۮ<���(�se�ϹMd�
+���#�X�{b��>'�y�.���������K����E$(��q���/�6%5Q��k�c�D�z��H`O��*g�CH����di��ͨ��	��9{�f�X��`���-�55�Za�0�d��x�o'^�s��ϯ�-Ͼ��X�:��Q���>,���8�JN)]�c�<�%���� �yf�iqw]�TC��5��L��CHvO�=�ZjS�VԐ�	��Ƣ��/�5;�S�����t���i�WB��Y����1(�$P�x/��� �Y�T��cz �$�����of*�%v�;�ߌ�yA��� ���%�ř��P�ה�yx]4�g <*��;����0�
��yk���m�+t�h�u�z�oZ�m��Ե�BR��ӄ7S���|x#�T��i�_������)�aE�s�`���J9<�癋���^8W��͉���5�এf\�o��aW5�\�[��S/��!*��w�ǼlmPoe���-]���I��cwU���Zb��l5�C�l�c��h�<ۮX$M����f���@��(�y��۩܍0�r���A�R�ۭyi��$D�qJ��g�u'4"�5�����<��������&��Z���M6%���`?�\�[�6q����Z�I���R�������#	y��6a�g0E��Y�LÆ
����� ��2���䨺�Y�:|��4��
�YĪ�"�-��N$�8u�"�r���^<8�U��$���"a�v�d���M�A
p���)n��~�)E� 0Z��Q�O��htw�dS�܇�F� Uۻ���`��#gӆ$�Н<"���L�M��Ej��Y6[����`B��&���~��j}�����g�BP�Ϭl)��Xn�QB��v�:>�@�bn�K�	��)v+��kݻT-��(�