XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��+=Z�p��Wײ�GM'�F2	���[�q�#��`���Z��Bi��)�S�Y<[�vd@� ^��1[8��5�ڸv��۶h攵�������#��&�D{ڷZ��IZ�ٲ�p��_c�ӕV�^�J��f~͕!=�������*�>� 
�H��SZ�3��B��$�����gs��o��%�o���A7r�=F��>�ӝ����B���K^�'|�l���`h�XG���asr"��8_�&�NF�-�Z��K�;�;_ś[���!0z�o[Se�$�ۓ��*�PCq~����*��jah)כd�����c53h��H=פ��m줎O�h&!aH����"�k�K
��Ѿ|f�u-�����3F�����=D���
���S$	��\���`C�3)�qޗ�͟/���,Yc�`�&��/�� :MG|����ٝJ���q}8�J�J*-2Z�o��V	����$��m)*Ru��7�Kz��y�q;��4��G-���T�l��6��� w�����K�_7��uI/�*��ň��&�m;�~~��P��e��C�x�Q���r��@.��v(+'v�i��$I������6�D�n{$vQ(��D&�$3����3 ��ܸ�4Q�2���:����,c�n�Rs��ݑ��$@�t{����s�@�x�x�'^��v8����<�&Oָ_��J��e8\�8y����u�{��T�VDvI~�w4/�U��
���Q̺�'�^lC�HXlxVHYEB    5fea    1830W
HT�&�DFS`(�K3��	KK��lg��AL�����p��;"�N�1����Z��� F~r�73��,��rw��<5����2�,����c,�)��cp��6��:i�Xa���ظ.��I�V�0�>���փT�F�{��`���<�a=��پ����k���u{���N�Y��+K�n Nf#(9����p:�� �a�O ����Z����S�s����%�m�ObH��DYԢfM��F�!Ҟ)����E'�� eu��P���t��W8�r4P�O!���j������%n����T���'�:�4�/`��+A��|P��*��5.���6${M��<��+�ŁO��k��Pq��W�L����Z��)B�3�N=�7SR<�-��ED�*��e�� �� ��W���ӷJÍ����N�%.P�\��:扄n�{V
g��G�4���Xb�M�*�4�#e�/�YO!��	�f�uG9a����7a��l4���	~�'�!	R�m���"R�Đ,0:}��>|����܃�]
E�G[bukv���-�zZ��'����5�{�г�:�R�6UFQNS	�n��i��hi��͠*�d;�[P���[�Ld�����Z��?	z�[�:o���)ҝG//v�Cw#�7٫XZ�.�Ň)���ɜ+��6�GtC�P����6Ѫ$t���M�?w�;'Re4�D�}s����?�c}=`�3/�5�Oߘq/u����.�$l�7@u��������{~����]��]R?k��K��]���\GE7h
a��D�	m<d�:�ƋN�{D2�a���o���+_��x����.+���7
{��&�H����H��!�!�0E�h�:&������B�[��v�=լm�8"�6�4�1�Uom��q�ܱ�� ՗�cYgc]����N5c���G"�j�ԡ��x5HH/�}s@~�n��YoO����2�Љh�R�-Z7
���2�=�@{�<��bSgL���_3r�yq��
;��;��(���/�Kj�Ұ�CXҜV�[]�v�
<�R��V6y@���<���>
�it
�؄_Z=X�ϗ-lӵI�DC�}�)_c{�TZh���ǻ�o/M�i�����X�+����7{��(5`�cڽzز�"���"w���'+7�*a/���5�C�`�fA�%2�ɵ���ʑ��5�6$L�o�Ǽ�̑9%��^��ؕ_�G*a�!�vw�8����i�R�P���S��
�`BI�[^D�~Pf��۠\��R/{!.�:%���K��v܀1�n�N=L�7NG�9��T�*�W2�%�S�^|�0���z��5�R�yl��$�lӐ��Օj�?)�k�K3�Xa2�p��!k�>O��:�J�#A ��������M�5k���ێ�:=�T�/������YŊ!����(���X���$$b��_����L��D D&���at�D� }�gɳҏV���q�����Ƕ������I�+�tǰ��Xq������:ӏ��qx'�^TP1FE�FI"i��ܹ$�ɰ-�כj'ʲ�a(��>xE^��|�W��D?�]?�#��/S8�L,�'� ���͒��'����t ��:=f�S~�<%.L/�n�'�o�@ ��z���{�?U�	@�z���~7�R�X���cQ��I��W�Q�����ak��O�C�u�-��PW���=J`�@�w�~R��TyMLϦ�e�I8�'H[��:�7��3���@d�Û_����r!h"Y�{1d{?�1����?m��06��_���i��8Y��H-������ՠםȬ���v�-�f7�C���n�G�ޖz�3	��y�?���d�I(tU g~B;7Ȣj$C�wk%�}�7��O�&黯�0@�]�vm��"d��RA�@7}�% ʲ�G`쁝R��qv4�W<$�^�te٣��3�;�qr�2�/�[jIx&&u��(����3�l�E�p�c���sK`�b���?�Y��N���l&��	�����(+�r_�$�J��9Az�+��c�����!������`r�R�e�)��3u��������%�� �q���mɍ�VR����,��z16��,���8F,����)қ�%J<o��V��#�.�.����h@��}|�}�-1�(k��5��m��<��,�X�X���3�zC�Us�`�ʫP%m4
#L��"vbb"�`�����I9����e\l�NĮ�v�t
�567R���(gb��������N��e�q���T�\}@�O$/��{��2r2�C�?��x���d��g��"��l���ct��?R��Շ�1U��	)��;�]�����9i����AM��nZF��^�XL����������a��W���Jó�& ��a�9��,�r���'
�r�UMw׉,�
���H�m�d�����%��o��IU~mPc����cj���w�.t���>i�fXS�&��Gw�
<�\̇��]N��J$N}�f"��ۺ�}��L��ޥ��H�Y+^;*`�k<��q�p�j8
9��������Xc��;�=z#g%[2vT�㥘�5k��l�aG�K*��������ԫۭ���5��s@��t����)K|oz0{&|���qM{��@���Ǒ�c�%���q�IV�� 0A�W;��MH�{)� ������d�����?1�o�&�qZadf=#<B�wb��lE&�Ӕ�1<f �Rn��K��N�\;v��~��f�wޑ����f����w�Nw캪�\����d�K0���f�����U vn p�m�Di� �p��,uq�E�J_�Ps��1$4�s%�%/W�Ӣs�������1��qY�P�U����8'��k��u'[�'鱹��-5���꺐�W�#� NQ�Hk�p\yF��u��@��H�R���l�
�Nglop���In��҃�?&�P�ZZ}����e�Ǧ4� E�X]�@�7L���B����v��Cw���Z=�,$�ˊ>��Td�8����Ӟ� �O CM����%�GTX�y�5��_��9\y� p�[_��<dڅ="۟���O�CiE>�L��s��K��|��<������g�U���HBU�c����n�mǫ����w��M��T��i=/s�U�B�?�t���1-<)!1�;�LLiX24N6�%���$�%*�@�J�ˑh�Mf%AZ�%�D���36�#bK�'>[}�?Q�y���_J��J�"�y�)$�z>Z�F�T�3_I9�8���E]U���)�}��8V��O�G��>Fsm��a�8M�`,3�r���e>�k����i"2�/��l�V6�S�3�����~�&�&�}�i�݂�}�c؍�m8%Ҡ�wrʫ�u[/K	�$.��Ā�	JMƞUAX��\�����.쪅mN���ۿRQy�.�����p^VF���O�}�x`��c�]z "��a�s�yuJ�_>%,�!4y�	��yD'�Ҡ%ċ����4����	1��� �h�������G����m'RHb����|q}���O�;i��$�5߼l�Xp���Z�C�����9 0}�Y�	8=�q0��8��+����㰭� �S��ʷ��l��L�E0
��ZN�5�Mw�ƲE/�I�d�[{���L�<�{Ѫ�J-�U�Ӏ|�B�4�Fn�9:��XM���8nR�a�t�ifQ�!�OOY��5r�27����������%Mx�Gr��F�8eh8�3:P����mW�Og9.i��[��D���~�2�Wi��H�GӦ���ku�iϖ�fl���*	������;�P{�ܔI�'�@H�8�3�a6����ɵF9&5�t,ev���4FR���h�S^�m~	1w}�֛*͸#�)��a�RI8���@́~A�ZeE��8�5j��~��S=l\�p���5Zq�K:�'/�������$t�`͔e���$�S_�1�7��zK/b��`���s��SE�\jD,Hݢ��>�D��E��7ޯN�����d����� �?\�i�|�΀��0K��0�h���5��@!g�Djk
emg�
��,HV~Ӊ����? �~N��	iG�RJ���6�����+B�_@�ո"�n:����O5�H���1:��*�Ј�V�Ao6�&2<��X�  �_�=���ն�pS�;��1��n��eF�?u.�d&���N�W ��3_e|��2�������^3ɬ�z _p7���h��2�p�]0g��(�~�dx��cþ�6(ArTg�i����7k
���b��SxM����j��g�}Ǻޏ�F	H�f�;�wR_5øz(��� �jB~6nt��5.ԛ���7&<����W�w7ay�Ky�
v�qꑞ<��_ �>FѾrY?`sW�����"�!�"��/�
3�z����P��Qֽ���+��TB;c�@����f\�^�ڎ��>�'O/V4a�g ��]^�p��d�9lK�m��>���[�e`���>]3�ܨ<Ҧ����$�`qh#L&a/>���+�)�:f�osWy����,��ĕ�E<�[h}�G�xW��l�H�@u��]��>Ӡ�D��󲀩$`H� m���]��t�G'#�{Y��J��U�%�H���7��C'ϓd��cT`:��ƣȬ��R"n��i��ɍ��@2upgr��峦�:��X��{!��n.��(K_�p�Wb�/R�3�6��F?̙vQ̝U��J���l��Ѱ�6?�S1���q��w�@|��ǵ�ԯ�Uc�Q/T�M�I~t�̭�)S �4����e)��ϙxW�|9��c��;>�
��>�v��C�_Y���CQuCi����܃ˬ�16�ڊ�K-������6�D�\<i����4����Pjc_�T���bi�ږ�^'�bڧ�Y�$�%k؀K1��[��e��L���dC����})�Ba��s�*��O|	Z�}�ԙMT}���v�گP�o�������*fb��e_�t��.J�E�C���:��j���!�%y֘nU�vh[���؁&}d�=:{�����Q� �a�	F�yT�2���d�R�6 ��Gʈ�����MG�j���o"�?FD$�2�*�>��(I9�DI�°p�&_������s��x��[�"ƅ%�ĴgD�ӖJ��c/�^[�pa����;򚊡�f��v�V�V>j�0�C<eoH5~\��W�v��s�7�$6�?�-o��Vu���0���w۵��S���缪t�g��(\�m��x[U�E�X��ԗ��F��7W��(\��T&��"�^�!��] �{>��]�4rǕ���:ca��[<g�r3���2�\��ƕ1����I�9�h�4�����	�;�~��7�?���Y(��n��@�����{u ��ذK�C�4]����E2��a�2	��Ty�(�RI��f.�Lu�n��Ȣ��v��D1������J��H���2�"�,�~�)U���~p8�1�6dˤ�cw׶x�nn{��}�s3ob���<���3�����V{�S���@�ޔ��i�m��s<|9;�����	�FjV	���%	��2���:���>�3IY�ŕ�O�@cA� 3`��βVй��J�x��t����{ٷ��2�W+����ʉ2�Oն�����A�[aS�� v�=����E����O��~�	~���ؤ�������h+*��\D<|vI�Yϥ �:���]X��;З>l�+2/�{���o}���ʏ����k��R��.1ԊS��ѕ|:��s�@�=E�\��C���|���Ҥa��غE}��(jN���le���W!��h>\�F=e1{pVKM�U��K��E�ӠK�ff/��Y��ʛNÍ&�YD��D.�%��7PF����,g��[�*�+��������]-zW�5YS�r[�� �:݅:vz��l^��������rl�?%��=���!�&)�Y��7�K
���3��"k1DZm�}L�G �g�R����R���0��$]�C]�/�	y�y�
a�_�eQ�=�� �g"���w�*�f��a9���e��M³*��S�3.h2���'�����dw��͵0.����!�