XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"\L�	�@�w7{��i�R4���j���s5�����^ޜv⦟�p�|���"��g�w��k'T���v���U�o����n��w�(>N4-��c0B�;���G|���̸����+'���0�V�K�P�V���un��|U���h����q��~\t������Q�t��λ70�VƧ�:����X�?����㋄֜��t��rF�����,����-R�D�J龾�m��g5!�p�;X쀎4�Y�tz�b�B�i_��	��.�7�:  ���\y�n{��JB��;z$��;m_��\�9�U���ԃ�\dV渟9�؊Ã�����Ս�[�[�GV�^�¶̟eu"���D�.��y��������s��u�kL�q�JDUǟ����J��C��ח|>n��r�T6!J�W��s��y"+	�ЗA����q�@KH蜒��ޗ�s�qjh���t�,m�U˩�&=��W�w����܅"S��\)����oxܷ���2E�iJ��VGTw��$u���ޣ��Q�����UP��X��o-N�1á�{o g��%���D�����y�	ym�yN�� }����Q�9�0�Sݍk&g(Z�t��	��rp�~Dv�f/�?"ƻܬ�m��!��Ȩ��Ǝ:�. ��VMϒ�cƟ+����9?���o�U��ؐ�O��;" ����'��o"W(���;��V{ .��a��������Vw�(׮ٖk[mܴXlxVHYEB     e07     680�Պ�~-��s��M᠔9V.>�0���j��ܾY��c��"�v>�����(�ǌ�^swI����;2A{M�T�}l��_��Ɏ�h�AT�ǁjqp
�������%���ԁj�]Q���RA���N���aȖf��~���"4�5�X���#
Б��~ο�m�	i�E/���LwtJ����z,��z'���.�W�֘�-�i4l�����|��]{��4 ��'#%�7@�"v8qCuB�A�m?K��̀e �	�@���� ��s��y�T830F� g�N���0�8W$JY�.�|W��|U
��܈Y����#��Ed�r�P.�jTĽ»KEy�g�Ye9�z򲒱�8����F{��ΚSN��`�p�]h�eL
���u��j���y����S�O?NH��"&qJ����m��- ҀL9��$R{����@}xձ���@B�c@�%�(z�<Zj��?�T'v��\3��w�2�H�����s�Q��%>e9��Г�����~G�N��<3.�W�[7;�%�D�G�*�m��1�����[�#e��u��C�ׂ)�n̑(*�Ib��VTr �1������ͅ:,kO���ZAm�A�g��EU�������SI���h��.��<&6�_��v��ƍ�[�����_8A|��C�F3��c�((�y�w,ϷS�1�Ky5�'OG�ԙ�-�WZq��H�� EpoI\�>թר���Q��E��I��'v�(ݻN�R9X�k!c��USnf?��jA���0�!<��2<܌���s!6���{74Wm0��x49RF�"'�±p�m�B�Rg�/-8}�Fc�d�V����������s8����ٌ	���7�\����a�K�p�b����~��
6�K��S��ۥ��j��[O+ �8L��Q��`���wD;wi�[�p6i���#��Iu�4&`�?}ʯ�xȀ�w,qX��+LW�"�� ��o�	6|`��Ia
��kS�z#�_�gh������ɣ"5ga:�MTv���Y]xAb+R��َpU�?W�g%#B:<(a�t��0&��6���2��ƩHu�����Bq^�S�/.m(>k��#�ט�{8�#�I%Pjҗ��R0l,�)l�vǮz���3ǵ�y؊5?��g�y�ޤ�K�j�8��{Iv�ڠ&�2%�O��J�y��1E���b�W����l�օ�8�q]��}B*
4�ſR�fR$�g���6�@y13�9����g^>��bX��\���ܜR� �zq(�V���Q!��]���.��`��'iP��;�)kd�m����o�ү9��.�Xp��Q��^��P�y�T�>�@���H��O��l��ת>�����̽����� ��W̋P�P������e�f()��e�$�����t��%#<,��D�.��Sv�^�_���b@������2e|J�]�\b	��F���	aj����?U�;��`ݬ�N��!����n(����y���<�H�qyI-�%�]2�W9���NPD=��B$�<�R?�~���#�ė��,�{�����ʛ�MK��%?�;��*],r$'\��BʸA#��TvEFBAPW�DN�����'Α4J2ܩ��Ap256�ύ�݌U��>