XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v4_s�$[C�e�dH'�]�44��۔�YP'��+M�g�ٍ~���U��Jws�wn4��Ljj�õ��T���s��T2� ;y��R�_��z�	��#^����X���esz�QYgwVJ2_����DE؁��`P��=?��Z,�OA��CZS:{N��5��qgد�!����kzyt\5jg[;���,�@�4�g~N�=*7���m��$���f����.,�@rJ�q���'M�����s� H|�C�'��2�o,x�T����F��X�t��[�|_�G���(	R�Ň�?�f|�+��Z����Y��?d�F{���H/�'�S�uK��H�����/[P�O~�b{�ʟ�l ��sb�!f#���-��k8��Ü;'{�t7�����[34��18w�A+lύ��w�_�v�#�ƿ	�h�g6�"��K��[)8�"ҏ��(8�HE�9^dej�ʧ=�)��Chv�lgI{�Fw�B���=��CV��{�b��b���{	��%�8u���Nf�6J9�p��>t�=P��X:�RH��!�qz���]��ޓ�>�.%��|B�24��\�#(1X$�Tz7H�Xp��ȅ�Kљ�u��*c������O簟O��i����:��ɮ������.��{y��TY��m�p���(tQ�5��jJx�KIL��ЈEH���
@؄��1<̃x��Hb�b����W�|��x�����I�J7�W��XR� ��z�BήN�mg��TU�D�Q�ZXlxVHYEB    95d3    18d0߆G�Mu7l(�+�f���އ������>����U%�d�lO��,����5ʭgV_��MP.�6��uQ��eR�m
d!�C��K���Y���~����	�Bp�(��9����:t����>B���#�| 0s;?�¡<�E��.����X�1�2rn7fi5�5�����~�4�2*2��(��m��BC�p�i��,��~qg_��7]����&o����\\66�?���u�5��G�R�!�G|D�-��3�V�p�
}�3 �°� ���	�/��?p���8U?Ok� �`̺��&'�siW�<�m����?�	��ׯ��o/�P�U�`��=��:T��`as���� �[�@��3�in���U����bs�$i�ȱ����{��vCԅKW�ś���Z��ŀ�}*U�^���~�'۪'%�r�#^c=9A/`pJaf�ݺ��:D�La�u_�5�Xϡ�B=�W��F�
>�v�I��e�c\�!>�i���:o��D��
i��-�v�Ҝ�ۋXFO"d���w�z�Zv��@@�'�vj_�w' 5J9�ź�)�^�a�\���-���al�ޙ�����ɓW`�-# -�Q�*A0��O�|{�^4u��a�`Ч�/C+@a>�_5m� �~���\h]���F��&��Q�,3����V�� +�(=o8�R����O��c��h��\���r%�i!���A�m�ھD�E��c)*�24�����W��W�~�<ų!��d�G�9��.J��'_J�ؤ���)�(��G��o2��ɲ�%~�t���&��rlYk�
�Vw�[]�
zc�u���<{l�+��Q�xP�a-���	�)�(2i.ty!2�k��4-|��#�.��c��>�KRh��M>G�f9AƽY5h� �z��*��{��V�a�{��}�/�Ynp7�R�)��s>ݐ J���)�| ��ƃ�e.!Є�DƸ��"o��YS�-�$Lcݑ*��!DG����I��i�42�oGL���6�ڣ�ߗ=�-��kd�5��|���A��@����.�;P�36�M�qQ�M��F�����5S�7@�ICi��d8��í9$���|��p��"���,����G�"��/����f˯�-��
M� ���tG�ID�s����O���m�LOjkh���y��sS�_�yzT�X'�����c�9E��w���͝:e����/�ig��:�C�뺪�>=]�@�)���R��=��� ������8�Hڵ��d�H���-���(TY|?�#��ձt&����m��#��U�
�hi�%I��fW�͞^��q?t�=n/�j�!a�Jg<F�)�	?ֺ���8�9��65��@��7�Rm�e��YA��/K��7U��jexl���̠�h9��]�j����&�����1{��rK�zv�s���>�>wj%5�VNɲ]T��8��I�vt_46��T��4Ѹ��Э�\����~ğ�2 ���e�1�>~��-����&`�Ym�m$�z�n�J��zTV��i�Q:�m�걞6L�S-�{�y����r���w�5���?���',���m��]��a?@�~�`B
��?2+�ȑ:kV8�Wȯ���k���0*�G�7׌M��ڰ]���|כ�pDy]5WC�h���q�^�;[)�T�g�Vi��w�>��^L@�Ɛ�ֱ	i��*R�c�dZ&�OKp������Vs�nO-x�7��˦��l�a`�T�uw+�����c�i/m�n ֿᆞ�59��ջ���my��$�I��*�x�~�� ��:�ԃ2�
%�H&�f�h��V����㜖w��ȣw�hW�&����5Z.3C�Da(�l�r���%A곆�)컄�Ͷ ��4�o�ŏ�fwB�\���Q1�c�-���3x��duKᷣ�YU[llc��>������	�δG����A�v��|X%���eY}����4��

�k�E6��'�`�?�e	�����>�$w���i�q��&����"aĄj�ˊǩ�y%r�XI���`kC\�d�9��ի���ȱ-~�Q�}
@Ұ^�p\Cc��{R�&֔�6�5	�SL����'qȘH&-���MO�3���Ux���R��Z
��gRo��o�Qi�饎?�X��X���,�w;�[������n-b#.�<�s�w
죚�1~x��<�������̭���9	�9Yl6�!	Q��8Be�K��|�c�3�����E��2&B��t�o\�3�7��yt�h���VN��B��ҕ������r�e�69F�F���0X�ht���y�JA$Z��H��t�̺{**P�.��Y&s��Oz�i����;��%fWU�עM��v�IX��nk��@���
Z,3�� ���P� �M���ˣG�?��N�%�^�_�Gn�!6I���C��uf7��Ͱ���n\z��jGa�v-��s�$��/D^��W������86@�BJ�_�V5�s��yjC�d������r�S��K4�1�ѥ,UH�y{5F/c��6�;����uj!��[+'*&��]�Cdu�U|��Í��ϟ�v��6�e0&�|��j|+l*ݸ�%�d|��;�O��K���ؖU��2Ev�P_w�ɺ��"'��}v�i�T�,]����� I5RC�����bo"n�u&焜�I�@wg�T+��0Bƾ�H&���
[�d� �E��>~��p�NPH�m�^�� J� U��U&���Nw�ʉ��±�Ad�\���ػ�:���5��~�՜�<���b,�����<�484�'��:������!_�%��M�K�x-�w����Ԯi�6���}��]����Ef��+�U���T�_��z��#<9��H�;J���G͔,GǇ�H�50E�K&/���-���Q��ٽ�#^=���[l5~|�v��W&�?��ls��|G��O��1��nz�K�>䫐��6LK���?�$c�״�J8���di6� �IB�$���}�����B�$�F���*��KE�h=�FS87��^�9Y����kb�[)����t\5�Q����hc��S��"@�DVY�L�\��C���#���G�5�>ܻ��2UJ��_z��oYهJi�b�/y�ja�K��}������+�2�	}��G�Qs��X)4�W��O������������[{�-���r���Kl������5Y�Yﲔ���z����������4��VХ\�a�^��kd3���k�w��|��]&�R�`�њ����.GN��~��Ԙ�T���'@0
.��O,�����N$~��[��N5���l��rr��?�ˠ�4��q��,T���+Z��az3"�O����dz��d�F�d����!�iT͞��:�⋵���\_��9q`=W����e�k�R�u��25�<c4񇼗����dWO�s\��I��g�LHs��G�2ݗ��wa���az;�%���9+�+X(G$��ԍNMD�mll��kv��T��%�gv�x��$?3�l^�{r����.`j@�jMA}&��M��Ì_�<�K+U%z��Kן-�B�9(�#ž����`��� �>ɮ
kэ�_�h��^*�����-]�Q.�o�ӄ�$���W�3�&����(}�:M�P(�."&>w��| }���	�=��(��-��<x���N��wbܓ����m2>��T������8�oA�9�IIe=+�Xj�H�H��r�5���<;C�To �0�S�B�j0��39�8��]��E^z��t.)p�=�;p~g��u�4[I�>Bɿ��������`v� �L��ղ/�n���|5vݬw4V@$f~�Dv
!�i�?|N=R^{����
���4U��a2���)�����P�-������)nc�nF��w��G�$�j~�7��\�ۢ^7�����E���f
�C���r8�@�')�,��^H�kz�w0�4	6��G�G�)�H����W��)g|���!����ͬ��ͯ ^�޵�v8�v��c�C���B�[/Vg�əƌ��	��P6�%E}��e�*5�U"��XA��M��|1�j��;K���t��F� 9�iHI��?$E��O��@�'|r�*�q��}1�`ߺn�&k)Z�ٟ�b-̾sj3ᆓ}q�bЊ�-�iP������Bl�NQ�qT�����1��㶲��ܡ��bב�`��+��5?NTc�����30a�d�v",�4$��b��2���H��!Ch,hx�M�1O$�Y:H�_m�)dF;��/-���+r�\�d�Y	�tmeמ���sS�ӌb�c��DN6R�r2��k�u�x�S�nP��)=���T���Ãm�X��Z������lL���Q�:�_��0q�J���ȸgD���|��W�ݺ���B%��T�5g���n���Fx�+~��&�#�W%F>���gU3� $]$�ٰ|'=�����m�"R=&�uqn��z��֦�օ�kl��/.s=� �7@Js�����MD������ ������8w)���R9���t��I��_��@Lǽqġ�_o�"*�{���3;bX��ip��{��c`�Ie
֪��}�"[J��D��?�b��W-fV6|݊z��Z�X)�AM�$�wϮ�5kJI,$��|4�Ѽ�7!,6����@�!螌�ܪ!�)K �w�ķ�'1�����f�ȳ<����.m�
"��j�5��4IZFW4J>i�"k��m�E�q�ڰ��z�Z�j��2J��q��yX=��~ٕG!Fs�?~�� E�r;�O�ƞ;����2��A�j!lv����Y�����V��Js��b��2]]mo�&�Ir���3�.���!$p>cj��|���N��ؠ������5I=���͵�����z�ݲ�Ø�+x����4?n���UJ�
|BX�!T�K� Ыu�l������U�"a�eL�~�zC^5�c��p�s+u��G�kBY ~&�Q�$�	��
�r	y�& IErO�V�0��z�NqZ�y�"^��O��{�%�����[�4UP1#�;������f��э�#���؍���;�Do�#��`t���;AH�p^8['c$R��O������D�-vh�AӜ����Z��U�-0�u//�=�.��!O�LF�������W-�|�]����&��Kx�#$�|�8����ӣ ����E����؆C����0�<���4���OS��/sS����o���K�7;�G<��K��w!��ԩ$���O�Q�C�4� iQu���n黷; }��%��|�ީ�:��}kz�N��F��9�Wyn�[��e���J�㻬(������#n9�=ҥs������#<�ԙ#�r	�;��6y��$�n��8A}l�v>�/��l����<cpЛ��>((=ċqw��r]5T��9�����(=�}���7�4gF#+���IB9l�j3M6]@-K��>����7	``�,���y�E�O*�#j�u�]�^��ܰ��IM�0̿�Vtt�����q�O4^���U+t���^����Lc�.����� t�=��,t��$��a��Ce���,�D��.���xL��C�@�VP+1��6/+c�j��(�a��X9���ɝ+�$�-�U�f���f���p�!Pr,��g�1���/���Ħ���H[r��n*y�n����]��g+�cSѨ�շ�{,��!�/��M����ѡK3�QZ�$� ��na)�������j1庞i Gx�ۦ������� ��ǮR^��/_�z`R!O�9�{pO{Z�{[6����������^�����/3G>��k��wuEJ4��L3/� ��f���F%+<��������՗���s�Hl�Z��$� ~ʄ�u����H4��������<y�!d)C�gH�{t8��Щ(Y��k6�Q��p���T��8�
���2#�	]��+9 �X��g�X��T9�� ���и&��߮���7p݇[&P!3����-��v!O��*�n!�~�I�����-I4R���&�J7
Q	� G�b;K'�ns��5+���a�(���a�c	�dfp.��]�*�����-���H�E�g��-��rM��ߌ�NQ>n�T��H*�n{�C����U���N��c�>�'����c��	W��eʂu��uRp�қ�