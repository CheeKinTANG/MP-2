XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��(�Ĥ%�X�삳T��U��?�B�(j�����l���mX��p,�(q���I�1�b� �C���d������xy��Z�A�:�i,tCtA�Y��ؼz����Ԥ��C����7?�2�(��p�8mI�%����X�Jw�8�9���ۏ����]��C;�֍��W+�!�� ����v$��+��r(�<'�@�%xY�J�u���%5��������9R�'a3˶4�ܷ�Te�7V�Ax :~�b;�qp�s��N�eܦ
�f�B猶T3y�~�8=��Og��5�9ģ|W`{�RV�O�=h�{�
܈��O�I������;�]`��Q�,�?����"�}zת��Bo�u�0U�<�E�M��F�[˷]U1�7B&e\�5U����CF$��f�a&=���ץ�`��zo�����d�W����T���d
N�@���rlA
�[��@.ߞp�B2�&����g�?�O�|�m��A�r�Gl;�<�tj@�����qB��32���t��Z���)s�Ug��F�W��Y��t7_	��A*O�V�vA}��x%tIb�;�\���t?/�;۔�����v5����|Q���Q1�G�~UP���C���9��Q�K6����A��\!�qV�1υ�6��"�1�?�B(���p� ���'n~�مU)V�fDE
{�|C�����!�t�[���~��#�23���~��J4ն�t� ������:��n�$ɞ'��1HF�]j�XlxVHYEB    fa00    2a40K-u�*3���p�X��-4
5�\�z3W�����/��z�`tt5$�7oŠV��]��yG{�z �CtKc[v���ל��8�%�4<�(��=撟���>�;w��4�d�ݽXB BB���0��\j�:t�f}���4cg=�UF$ˣ���9;��$�i�DCU$�E��ܺ0A���K~�ɼ?��y���j�#!sK.�ƋT1��~�Hנ�Tf`������7;"���L)���
|��KP�
/�3R%�U�8�!5����E�:K�#�oR'���������)����_�˞,(B�����i8�Y���h���\��)��� =�>N�Val��-{((��&M6S(��JyD����L4!�Z���E�g���{i�s���zg�!��T��4��X��Eg?��Q�]���� ��:&u���"F 2���$�oNѱT��ЅO��| C_��^��z��vn��=����u���<\x���7'R%)"1��m� >1��B�zԍ2�B*�]Pr&�ߧ1�.�5��..�{^@Ҫ,w����I}�#mެX�(a��>���q9q�N�[9�Q����I��'���6ځ�]3�O�Pf�غһ�`Oh�RQ{�����z��L/Թp����fz�@jQ��cۺH���|.M�J8�ր͇�o@rA����#��w���%h�����p���&� � "�#r$F�� �Z�fξ�{IH`����x~9���Ȟ��`�k��]w�:)�؈n��C"�7d���e���������±��;Wz1� �!�@n��Ԯ&����� ��>{�wҀ�/쐧�µhae턅����T�T.�_>Ke�BϢ�*�/W�7�t6y�Ȭ�]����)�O}��T���߀��ck��^���֕M��]���;wLa;0�?�rʁ~=q�<�L���(��h-�����g8���U�Ϩ'��UL8�Xa��C{�!� L�ԶO ���7��m�a �1�K�6ys�܌�
����dJ��Р�#��D1���ݳ�;�j�ɸYt�8 @ξ�?��~g��y假F~�*��L��1@�%�G�`5��$`��aȀW��ǝlD5�K���%B���vhg)헯ҽ��E�î�VT�:Hq�(#�t̋�AeL##*�ڸI�s��}�Y�M�{=Q�4��svM�5g�vt�~$x-�P8�h����/9��m��D��i6:coBI�O]��`�[���C��S)O��Npt�0̫Z��g��P
\߮�>�6�9t��[x��;+Ua���r׎7�ɋ?Pw���0�c�Z�4n��*t���p�.K��Ӣd��Y�`�Ϯ�D���v�E�6^<!��6��Ѐ#q��m�e��AT���!�c�6���r^hX���a]�Oh�P�`�f��:KM������տ�3�!L�b�QK�q\Y���)�Ue��Qc|��~�v,��Ed ,��0��U��Q��pB�����'RZ%ukźm&��0��#��������F.&*Ɣg�?j�!oR��ɉ���w#��?t���c� �rtG���xր|Q���>Eq~g��鉅�q�Kތ̺:�#�L0�NYJ�d�$�*�j�� �$<��O49�-U�#�A�Q;�-l�*pM�)���#{�RDz��Q��\�W�eLYʯg2"<ˈ��3}� -�Ax�=�e��>W�܉;�ńsX��]��ڙ�F3j���TM�o]�F�ej�7���q� Jɩ�6w&��Q�2=.e��F^�:�#T����5�v�M�jg�����I����&������WL����oR#��?cS���$w"Aܢ����;�O����c?K�W/ɵRD�U%V_my:V�CR��,��͒I��Q�!�g��^<�d�_�~%SVe��=�J�ԅ{W\@�%�-s;�s��`e���%��}`�H�T�5�!�)��q��S��aQ���0q�!��q�(��VWPM��B�O�nc�>v�x�J�����p[����?}P�Nރ�]c�r���U@y�b�a�X=z��L�e��ժ��c,�j����T�VX��%҉��ߝf�Z�|�r/`�J����5M�e�Jz�j3�U[>\cscn�Ź�A�y�{';��HF����k~�����;�x�s���@[���j?�沉_��q�'>BN�ȫ���D�jy��4 �\�n�x'��j}XhO]�j�]Tֆ&m�#?C��H�<�A[Thw(0�o:X�$K� ���-�����g8(}�4�	qv"BO�<���h���Z�)]�5�3���zaŖTt���N�(�
j<.�d*��䈒+�P=B���K�q��h��}�Ra�3���&�3�Ig%�����`����?h_L�8Y�#���ul�9S��I��Yf�>R��g�Na�<U��IPa:��9��{+�u�pC��j��1�����wS�Q-R����>��f�����c�)����,�� X"o"�"E3�U ���8�>�om(	"<�^Q|c2��3yWc��;9�Z������	�w�f��-Q��G|�4L��%)��3�cY�-2�� ���#Y��4�C�G\����&����߬�"@�Ǆ��\�Q"��P��\� ۃ��v��e- ��K~G���A��oVq��,:�wVW���*��u_��J��Iy���T�Dy��l�(z���y��߂0sy�Ze}|$���H�]�qG�ġ��~�/������z�+�>Gb�~�|�c�}ܳɪ8}�	x�tU��胒������S�e$BK|D+��� ��l�FS��yD��M���x���s�!MC���O����5ᙀg�j�Q�����g�����fU3��\����h�i�����Co�T_�{L3�f"�ߑ"��?���ߥ�H��9���)V �^q�i���,���
�����4�,{5���@|��hVg��Պm�=驟M/�W��c}��R��̒N�/���ϢR�=�`���6^+k�x�̢_{��i���1���;vz�QFZ5+��[�����5
t��w��ާSj�4	������7�����@�M	�%*�p�*��H��~���0��^�Y���B�@����Qmfa��h����
X�n�T�,�M�������W,g��-p��_��}.�?q�-��׾̃\w���6jJ1����2�],Ȇa�A�Q����|wA�an G�F�j>��c�/��S�bT������L߃g�u�:�H+)�m�Dk��BsrT�"{6�q�*d�ST���l�?;���.��
�e/R��+�3�������8�)ڧ��A���Һ'�f�z��~��e����y7c	���S���-��������}�u����cH{�Px��)�]]���;}O	O.u]W�׃��f��na��5aZ|��1�+�ka�����u��r!|~�!�4�4Y�~	w^Y800u$d7�O��yE5��!������R��K�+��+�e���?t��i9�g��u�js�?����vr:�!۠f��3��?��_`Ƅ	c���qS��Hqc�+�NX���nOz�s�v
�Y���~
���b��V�Ԥ$�T�������p!��g>�^ �裮N��1z�]�w�]|�bRq��n��s���z-עq{L�������ywB���I�TWB��/�v#��P���p2`�1Do�����jo�8aı��m�i��3�G�pس�l
� �A\�c�$ �?ՇG2JR��F-����?�q�i��>+3��XWkd�˛���m�@d�-����&�1Q��Z��BQ+��)��P�jD2����ֱ�h��n�t�e-�#�RN�iT�� �4H��6x�r�rFR�-�&�����d�h�.��g��	���{L*K��?�K�R0���D��¼vt;X���J��]T!�Q��]&b������S(���ɯ�A�����k0�dB��1�p�ܥLa�	�H͌�'�KC�VG��idP;����%����T�/tS�����R0���I�p�me� ���F����o��qŅ�`�p���9@m�PJ{������ )w$�j�+��l�
^4�~��46x���@��񖡞]�=<fU�p�c'��]�k����m�ݢ�rޮ����P�}�9�1s���Xm�ը.���v�RC_4 �c�7�s�8��n'�Tz�����X�c����n(i�^���l�y���A�("`���؜8�LPSf�Bށ˙�K��X��5}�����ĩ�v4�x���U��.!< ��Kl�Z��s^�)#�C����Bq��<��9�UwI_̍�p���g����c\?EqN����Ҫ��(��>���i���i��Q7���e�U{2U��,ϫ�6��C�ľ3�RGa��O�S�f&[Ft��$���F��;����']�¹��ZF(<$=aÛ�z?q4S4$�W����M���Rj�6���Ɍ7d[�%�I�O�n�L�a�,�k� N��<�]�8#^F��S2W���lVH����O7�$-T���j-A���a��K��i�W'�`9�/va�~�Wx�\hLmL�g�o�q�V�����H�|�KDo��ހ��:�&:^녳P��2R\}ګ��HӾ?V�����pp�B�o6H�o����6�?�Ep
���fī�QG�R]�� �ƻ�����oQ":����$�@ɶ�>3C����s���0��[s��"���'�����XF�2s�*2s�0��؍O�Ky���gzm��i
1��H��� �v>L�n^O\��76��С�b����jҴ�� �iH��!�̆�b��gC��)�|����#H��<͖ڙ���ˢ�=�G/��Ke`�'۞A�ȁ�.&= M��(�6X��EITd^�N�Ys�O�@6Y�T��2-�\�/政�J�pj�em*2���rL��pz�z�A�J�w:��E��ļ���� �n�6l����?d�$b�#ZZ�rr����Gn=�����D�t����ԟ��ZѲ���pk�#Cf����V��P{6�i�'kݎ�Z�<p9[��s���Մ)`�k��u��9��_r�� �~�'W��S�7CU���s��* V$�z:����m�ܷjX��ikOn��
wC�2<�k¾H?�F:58��H�R�r���W�Ό)����0��c�������PdQz��|Ҁ�����+�c�K���N��H�����}���;1m*��I��lZ1����N#����p��k��+Ng�ݤ�\���fw_X��'NB���^C���22a���y�K�hb����U�@bi 1N���>�Ssu?[�����25��a�P��.�g�૗�MS�W��f�iPX��|�ΐ�:�� ͗K�e�l[����؁#��O[�Ӫ�-X<��$k5_>|�0ç)C�|��?X�݀�k�k�m���!0T�e4�
���P|Lr�΃�W54�y���ˉ�>�-89{���!����,��n�]]iz��hĜ t����A��C8W"�ǝm�SS9DA+�월~u���z��~����	��!6hK=�5�S]�r�at�Jxɨ��N �'��Ή7�\�*�� �O@��u�$#��'&RT.�%�ŉE�UJCk^��`��j�¿�+��s�rf#pg��N�u��dEE�0t�vMr/@�(�0�����=�x��<&Z����"�P���k5��z������K%lrn���n��b����o_g�@qyīߠI�Ѓ{�W���![�IDK�0�'v'ՙ��J�U%O|Ԗ���EaT�Vpe-�y:*�vc�����D��^P�,yW�R��I#�s�&`V�������Nm�t͍2�����Pxq�`�Q�46�:�Z�ZOy�G��s{���Ll���[�h�\����Aw�	�N�ø3��NJW����Ϊ�(�#c_�ف����ҝ���z	_��u�<L�7�ڞ�&2��o{���[�O�9Sq����J^�g4}��I.\H8A*�5,At�:��ӿ}�דw��q��`8�n*��,�8�6�=]Yq_T�[Ķ»��q����'ώ&����n�I��p�N�����>0#:?����[���Y�u���K5�I:N���|qN�kT�����2��DTm���Z��"��[�Qf�c$n��m��qk
�Ah�����X�A��gG� �Y���P��s F<Qw}9�	>\�r���S�b\7���J$��_r��B?%+�f��H��З6p���	&{~(X�AE4^�R����� Q�C����q���u� �&C-!������qZ$�2C������4��=��8E1���1���b��5��R�!�`N���v�Kj�����l� t��g6U��L�fM���l�U�ՎX��1��m�0��L������Ŀ����������+0@� 'u��?G��ՠj<����uA��3�y��$��g�X1�
N������5f�sB�����B��@gOC��x�|d��Z%��Ա��W&0k�M�߆�6%���qq��o�T��o���mS�T����,5����|�?7�^�H�=�qn;���[������%��Q�%7�l7�k�a���QpjY�k�Ec��٭@��Cz��	=h��y$6����v��yV�@iNk��ĳ��C�H5�p�-�oUv���ޮ���o>�N-�k�\􄅲G��!�Cꪟ	8�hs#�����b�_4#���\۪��=+=x��%n=�V�]W���־���\z�E@�6�g�!ݴ��<�?u���`.ݫ�on㊅��ssߎ���d�0��<�\���tY�>2��$�����h�����-����M�H��7�Qv������u?m)�zT�$ʹB9MQ�
�/'��>ʵ� ���Y��bb�!W�����u�N'����"V�t�#>&ƅ��qOnL�荚Sʕ�PzO*��4
�>A��|�8��nD��)���;}/A����` ���B�R-����{8�C+��c��O��4�������x�PTF<�~ͶD�XC@tn�Ld��MF|Z�Eg܆;CF���1K�	�<��@#v~�w����^�)/���m2���:�~a�?�κ�"��G<�
�U~�!��ʄs��Kv,�k���^?�خ��z���T�z�@����K��C�$�j��|��%�^=e�Ѷ��g�v� 3y��S��k���P +iN�6*�x72O'k��l���h�t�Ll�����	�AеͬJ�A$A�t�՜��_���AA� 0��<'f��B�<����}�/��O�y��Ť
�~��qҀ��P��� M��E,��aP��o�׫�8�Ǵ��@zA�q�.��I�&O{cq��"Q�"i�k�(#x��n�'���A���A�X1bZ��Dt�A|��6Om�7�ŉ�J�Oc��#d[/-���!~���p� Ê�Qp��p��2�c<����� �u�L�I����S��"������iB1��-�-xYb<��� 3�΁�G����o��E����+D��B�Ħ^�p��0[����V��m���u�j�*���Yi�����Qu v��� �K8�a���ta*�k"�������v�HY A�Aa	B}-� 笰=!�p���Հ����{q�������v�K,��M��,@A��`�)�&P�1@[��t��J��&8�u�II�YE���C���Z�\Q0���m/�&	r9<�ÔP�$&>������+�$��������D���6�Ge��j^�;��Ti8�"� �ԐK7�ʸ}(⍸[�\8�Ne�t�Ӵ@v�Hr�i 6ծ$]��L�����)������I�������n革�<�(�a���l��*�H��0��$A����dw��.ҿ�\���E#�N	���I�1ݭ���]�4,��a�ԇ�EmWKja���Hz�+z�23�F#��������-�8f�iR9�s�r�����.%xZ����u�/5�+,�Bｌ��J�	�>{5���^��8:y�"KE�'൧rx�	s?�zj�߈أNh�vmvk�柙�R�w�U�9$Sf����0���=$��k�N�~ʃq�i��b@@����ڎ98?��I�����S�Fܙu��9���œ@���vC�� ZʕrWg�'�SB�6��&�qp���j|�<]�����Z�(]��`�^d�8I�w�Ɋ�G]����Cj�G��]��p�Ƹ?�vD��k�#���ܛ�@O��)o�R[��E�ҟy�ݏ;����2�SC��y��E	�/�H���d�?,竦z�Qx׹~M"X	�Ms f:q��۫j�!�����SY���m�Bk�8҆eJ��"�,��ۇ�a�w�.���r<ϡ�y�	Ћ��G��y*<��o�avٖya��"4c���h+�5ʛJ����Qw$|��lt�Vvꊤ�'_�y�-�5gT�L��C��6��ݻ�N�T8D1��+���Y�3���Ӏ���[�d&Ǚ�	8z���t���2���ٶ�p��3qff,®�.�k�������>�R]�dOQ�a3�����A랛ը͓u�J�}�vj\��҉�e��QeO6j�y�8���{Z�8�oCՇ��t#��-���|�|��- �u���8���7�X�i?:�?��B4���ξ�}
q��V�}BZ�rN�<�Lبe���f�6��N�B�����D�X�B�^D@Z˻/����v�&�$j�Ĵ��j�Q�*(���WcZw�H�f�dd�ѝHh|c�4��o�I{`��2xr��p�ܾ@C�w��/բ���Q�>"b������s{d8dR0yF�w�O���R{ܪ��Y�~��
��k���D"��?����G���:��˰���ǒO��Ô:��'�S���}�K�࢟�
�����g��"���0Vw���{Co�WlXv������ g�\��we՟�.���;��r�ؚe>�5���QmyK��?�|(�a6�
Ǡ�F�I��U�\D��	���0*WW0Z�.-��Rֆ:����|#i�6i�!w�����A����M]�~��S�9bԤ��6�v�τ�ho�Ɩ,�kyj��Pe�4�~5^�����x /nͲX	͝�BC�i4n3��b_�}=}�y��c�h��.4���B�#� Z�%>�F[��~v�i��a��b�\�N�&~�O����a��!סa!��Z	e��S���C��4�`X�5�i�/h2?=����=s�(15�x@�g�;P&�3Q�nN���$-�[�m����)u��g�+b8���ԂH��?;�)
b|�2��,��J������73�{�Q#K��j�5�Zf� �4�����祚���Q"��؆���~��	3Ţˑ$5���щ��^�5��}ɛN�Tuzd�`�F�� �/զ)b0�r"�ۙE�L�����j������ˇeS��e��5�nF݈Y�}�RK](r�@��.0�]5��8N�}�~>_���J場Q�<���LT[��Vq�6�q��6��Ǉ����҅��;	ΑiK$��x@ ���:Jj��!������tt�9~B��`�z�W�� D?����ȫ�K����\�!0Qk�1�-4�������=���"�UT�n/�T�`h����I@,ı��K����G��wR7��ڶO �:O�̎��5��c�h�D.�� +�!ݩ~��y6��})�҈A0�7�:N�Q,���5W�]>{u�+L����pֺB�=�"bjTj�5	C|VNR[M0tUV������cc6g��	)�TX�E�����@��wN�hNѾ�!Z�e��{�u��.�n���QG���&
<m��k,���=�u+���(���9)��Y��.j�d-�l Y:�ߗ�fX�*}%+������ߴ�_Ab�J��g�ɮ?�"l�k���`#&�Ӕ�9�h8,�0nqv9~5F�:p��
�5����.Z����Cl�Nu�Apg�䌶W�@-"K܃\W�}3S<5�s���R.�|�
�$�Ƥ�
K
���o�F	rʏ0�5@�|G�\Jg�,��B����LAq:=�{k�W�� WJ��aO�`p4G�,�^��64e��*4]�@+�D�-���R7)�j@hHA��L�bS�?�~�Z�[\!R�('��^^ФLE�߶Ԙv[��IdSK����>8t/'f&�L�Ay�o�v~����Ў;Ϣ�6��*�Dc<�fC���=�(w;&RV�9} ?"
6"z�{�u5�������AT4�7{- 8�>�'�Uh��vG��:i�iW.��j�h�9b�����m���	7~>���L�p��o@Sņ�	��K+�&Q,K qsV<d��O����=��E!��X���܁f�p�����B�bNJZe�+	W.2lM���WEO�2SFL���U;RfP.;�qVY�o/ɠ�e�
��9���w�6x}P�3;�p�X2qa:Dq@�~�b���([qC�M�����a��w��NЀ2�Q��Ѻ`��I^�̶��:��|��9~Ak�	�ف*5WS N.��µ\����Ŭ �gI��"�NS݊Y��Z�4
^qB&ivf����\yu\��X ���meXlxVHYEB    fa00     8e0!�� �b�ZW5m�k��}܅�Y^�Z���#Yd.�m���n�����,�m~��(v��2iutt~��F1��V�d�#_n�y�c�}�ϸ�E�kc���^�#2����&�VT�.w��G�r�<��q�bM_��ގ|(�@��p}�|���v��=<z=���c���� _/��v�tc��+&�/?���ټ��l�b�l`�_�^������߆�� ����#�DY�@M�=5�t�c�������}��idJ�i)�6Gp�j�����T"�c)�?hu;�Ճ�6ғz��N`)�;t��]{��'�j~�݀"$�!�n��nS�I��x�~?��%s�3 Ҹ7����D2L�ä�+� Ta8)y
!������;{���e����M��O�9F����{���ͤƒQa����I�}'O������@����W��m5
d ��ut7�.҃��ӕz�gS4�(�z��Z��d�,�O��9�ި�yp��mƭQ�K�:ا�t�0��>'v��ۓI���Ϲ������cA���V���a�Uv�e��u�ŋ�A<��Tv�R��(�?$��'�盻, ��t��f��n_(�~0���>fb�@"�	-��	�wm�E��'��;�:�Z�M�[�G#�X�ϥ=*�S�h�NwF�8ȩ��DIo�P�h�]�F#sF�=� T�!�.F1�hj
ڻ����z	�Նe�;C��}^ɥb](X�y��'�W2�\�+���gs3�L���Yv�����	�+�_=zt[���~�w��ݗ�����_$�7�b�hՕ3��4nt�q���KS.x���W�=:��s�*�ɉ�2��\<p] Il��Xmv�s�=����K���j;t���N!&E
���,���{�!h<��߻�v��=�S9ȨDN��O	1 ��I�=7�)Ӝ�]�q���P6��i)4��iųd�fR���4�Sn�� ��	�W�-`~`9Iì�J�P�|K[A4�m�o+`�Tw3�i߃u��d�y)i��w�\,�r�ņ���'5�PxZ}�/�2�����l���˖:��eq\ܲ�LB;�N�@��p�{C�����X%����G�$k�Ow���^8U|p�7�I(@>��:v��`E!� O����*N�Xm9� @�	�~p�%�c��^��2BNOf?��~+�z�@a1{et3
r��kc�\��Eɸ�7p��̾�<抩�z�c�P<�����t��+��z�h�����H�ry�=�HK�m.��9�ť*�O�?������1�t���P�PЅ�ʴ�<0ATPW�(2���R����W��0N�fP�T�~���[�(�K9>9��$Ó*1�`Lu�rV>h{Q�[��ph�k_�m�|l*QX�u�:�9�i���Ϲ4C	��ŭ���0�\&3d���c���\X0=��J�oc�ו��U���Sݜ�[MS����0�(z���|�"9���[��9^���*yYh�:�J�Y��i	ْ��1�x��G
���W�"�V=8�5j?gcdLX�������̳�S�9�]i>t-i����a�s&#��m��/�L�׋U���i��3Loܒ+&���)=����P�b}�f%�s�b��?B�Y;L�E�o��ǀl[	`X*�r�N�eh�y8v�[�a�`���p�?	�t2j�8w�� !k��	��@�+Tj%�v�,@��Q��ə
��b,&i#'����j��%�5�n����	��k�V+�fL"�W���e$ }�b��-�,+W���☋��#�����z�HJ{������[Nq5U��_��eA�br哓J�+���N���hJ��8�rn=dgG%v'�ʆ�G�� ���w�U^��������^�%����ҪG�pM�w�Ԑf��R	i��>�=�� ���.�	��}2�7C�LF�f�n���sj�z*���J������0�X����۽N���wqX5�+$�'�ǖ�ws��Y��\
��c��盧�tāu;��o�P�ӫ;����)��4V7�$�n48p�%.��*>.&gJ��i0�g`��Mݶ����~<�A�!��}�]*��36
�M�0�3`Rr��Tv3%�xh�P޿�P\b�f��,�5�SJ�jM���#W���U��29�0�5a���〫P.!�k쥟a&�"啍�\ղ���D��8F�NxG�D��k�*M)�1�s0�z@�c�Z"jXlxVHYEB    fa00    1110� �P~����g��hw 3m��JVq���x����Xu�[ܟ=}��!q��L��߿h�ys���J�_-��a�Y�p��'�W(�MkE{C��	l���~�O������Ϲkjl�����`�����;|s������*�����ʺ��05����YVrb8����dy'iveۏv���6��ڨ'�y����̖�2�ZF�o"��ݜ��8|��,D�yj2�gh*�^��1��Ur�b8����\���_���.��l�� ���8���,ṧ�x�d�U`C�y�&Ͱ)����6��r�����������AW7qw�5�o��\7L4�e�4�8�l�R��@s3I(���T͜���M8�wK�%���~��_U��V�RRP�>���~̉�Z��T��`��k]Qk�:�\���|0s@+�w1_y^m�D<!�o�U"�8"��M��y�~��q��;L]�~�h�zk�u'~Bǚ�.�R��i�ڤxF9�ͫ���� ��t�s�an�8��g�F�j-�I1��i�7���ÇH�z!4�X�J���/]X����
+�/�'AY�T��6���������Zh�1+��E�ˑ.���Ȏ#���	r!�f�N�Yi�p����R�|�cۛ�|)�i�z-"�W���Tnҥ�R6"f��7顆;����8��{%u�@��q�ؼ��pEI�?͗����Wg�b��R���8��௞�l�8��h�ʢ�:��թZ��!��R��r���Q��r�8	�/:��^ܧKZ~Z�hڕiCѝG:��;���iF��L��5'+y'�bP���&�$T[�D�?n%'h=y�[���_���K��>d|����4���㸊�l5����v;�	��M�{<N������xɐ�\�/�j���������z!O� @LZKS���*���J��(q�*�4�y@@`XM�ys%*�F��i~�X���]��x�I���pD>����	�&��������_1�hu_@��Z�&�/�}�M<���h6���垩��iZZ�g2��~WX���Ry��X*�"�ҍ7�����y&���#3jS���2i���^죟��I�c��~G����	X�4�@4���(�n��+eK
t�6�X�bb\�p���WY�+%[���\�@������du�_�I�E�$��0�2���<`��2��cY�#L�;���`�������/��:����WЅ��ЙI�K��'�7��x�����zPx��+�I�bMNK�YyzV�$wu�5^�5^2��qI��=��T_��:Bqۅ�?����t2��@[�`;��8���9+_b�3GB����89	���|�\����&��@�<�N�iI�J�G���,*E��ME�z3�LX+�o���,����#&�nզ��>�ծ�x�jB�ǜ�X�hW�R�Yu����rx�J1�g�]�v���b/邥���Q��|n��D��+5��g����=�-�-d�-σ������Z1��Nh��
g�1*h��̫��:V�����v5Pz�s ��)��q��R&^�d����`
�������%���c�� �!�<S�1ñM��: {c�6M�+5ʹ�>qJ���cBq�W��Z���I��n�����~�ڂ�'�~�����.��_U�b)x�(N矂�a.�NeS|V�zi��^��_����ҽ�Ɇj�&�B;wp�&�ekz��^?[��Y�j�#Ÿ�2.*�,0-�Y��˥�a r{Μ�Q���F�6�3����_������2��:���4��	�56Uv�ށ�_ΰ�e/����j<���B�v<�����L貪Tut�b���L,�*�e�!���AmF��M��p��85}���`q0���9')r�)#�S[�}b����&�,懅�:���?�]��w��RV�e�2i�5��ZhX�T��v��2l�[�OO��&�"��	����*2���7�x��o��>w���5'cf�#�&6���IO��2� �۽�x��mq�VJ���/�i�H�E`��O$K��4l9
�4Ӹa8oq�x6}�YuY��f�D��^-␃�qr�k��x�����ur�!J�:������w��F��/�M՜x�7fK���h=����g'�.��z��+�� Y�xi��o���W�}���ő�>l!��W���	>2�C3��)dm�ta����g aj���@qAm�>k�|�"ϙC��̑8�&nz�� ���̊@[u	�	�צ���LI�\��䎒�]ed�B���Ic������!^��x�%��q�<@u��s�)MU�TVF)�� ��d/��ɗ��EU�䠾Z�[y���[�6�z0�\ۮ����gR}!űO�b�M�CT��9�N%L '�H*�OGdJw���	W��4�l"	�s�3e��gF0�>A�E�
�(G�����_ϕ3ܕi�\��?�(5p����5J����������B�*E��>�묦a}-[�d��O,/=�[��F��*3�B�GXТM�L�{m{�rM����u �ʎ`t�TZ��rl�3�3vvQ�h3[gǆ覭��8m�"k���u�ڛ�Su�i�qƏJ�������9BB]����E�M��%�y�:��g�v�j=K�MFTM�i�[���Ÿ������V���p�`Y�4^�Ui��GD�or���@�[���ޏ��Tm�v�Q�$e�Ǫ���΁M�}�)i��x+�H�J��2& c�S��R���8#k���K)��Ò�F�W�f�f��z���1�a3��J��rw�굄ǯ5s䦞H�.])1�ޝ-ٹ,z?��ՔpS�\LX��(���c�:𰖬J���Y+
�t�E��x�ų��㛷���S!s�Kk�dRǖ@/��\R��<ݟ?��s)$��-2�Ҙ�-*
��'�{?I%���_��0�I9W���o��4��j��0^������!o��y�-1i��.3A�p76����'�I��{y���4@��3���v�	�p��<��!n� Fó65_�u2��T�!�����D�E�E����~�o����,T��uɶUA�h�Mz�;-��"z�?vD�'�E�q�)�;��;�ϡÏ�!�I���\]G5M�fė@�"58�7��^)��J�D{��ؼ��ߪ$Vx*�;V�%VW�
�y'�	Q��B��܋�i=5��s�Bb\�OO	ax��3}�u�B8�U�`��է�?G��(�;2�v2��x��b`����������V�ʭ�.���9�^Ǚ���#g:�^�r��{��}����bfd��y�z��y�/��0�'���J�w�M6�o��v�#Y�%g��]�h,�A�Zx^C�"�yWz���rg4��5 �h˱Hmz"��K��ϓ���vM3�~�����P&�m7���#�|���m!��`��B�Wu?P�-j�G��|nF*��uYS�
�-g��Eoe�.Nqي���@R��O=���l�ĈJ�sQY쏚�/��@s��)I��C#(c���"�
R�%��>)�,�â�5�@8�77�l�t�dy�lb㟫)�%��ؓMi�bv� e��̷H&��2Eq,��Ů2Yrб1=5�)����^��x�S�Y�N�Q�N?dM��2��<��"7uW�Kјz����Y��}2���W�9a��R~�h�7/z�K2y:���Kf�ҁ�0�8�9�mc?U#+�HůZ�HB��%�$H4?�j [��5�`���wͮם���R�֕m�n���ߔ,���5"�摓U]"Z�k��;����߿'�P�8���@tC;����p6�$�W5�2��sƭ�����>�i�~�"6�l���r�c\����m����5�	��,)#(�P�?�q<�\^�#�w�ZY�Y$?SȑV�w�5�u0�M��BlO8�8����׀c�i�BtSY���q̿U�n)�#��?���|s�����y�9m��s�@f~��L�@��c�e�x��:���t�'�~`kg���d:�Hb~vV�eR���=�9=�F��Z2IN%{�������a�wV�D#ɫ�r ��In���0�xi|i�L�oWٰ�_�M�g*x�<oY�_PKD�0r���/u����NJ���B����ƺp�,-\�t���c���@�8
����JtJ���h�Nn�
�j;H�� ޸t���3,�)W}{�~��߭?�C�u]R���z5I��du;=�^��t�~�d�1�'��h
���n֦�E*+������Z>��qH�e��"����uk�#"�NW��Q>�%A�F�H���C��\qw�����_�$�ǋúXlxVHYEB    fa00     ca0-��\׵��ɤ>)�W����o�(s)�"�⏘�%�9W�r)�D�����H��m�o���|�T�h�����-P�-,j�#�!��=��<�|�d���H����;t'�K_Sn-���\��v0�&g��!x!>����.��8`d�E�v�^pw�=
��;���h	��=�������8ʠc@�c\���Jj$v�m೏��Fccۇ<�D�ݞ�R����^h_�{��O�b�W�E�Щ���}��@r�nqy��L��ܲ;ߜ,[,c��/�y� �A�а�OV��~��"hl�JP��Qs��c�ZdY�w/�ܾ����e�5�VfX�O;����uo�}��D��؈<�&��̌���H� ƒ����a��xK��׫S>q��oR�&�~_�{�"���3ba���*����y���y��#~ź�� ��xd�5��eC=��y�P��Xz27��JY{��[gɌ]��$3.5=��qM�����}�\Ţ�x L!}]�e���k�a�"5w��M�t��~�^R4�N���͇�= >���6���'��f��'�N���b��ҫ���L�%�}֧�WZ����HZVn.�4� ��6����Ҧ$��@U]< [�K�o.�B�K��H�vg��V�3�]�v�u
6P�]Y*垇?A��|������M/St��:��ʏM ~6��],�,��`.�o�2I��8�ۆ,͡��4Pܱ�m{1�m̂�~e�IG�z��p{F�@g+�t'��8-�#�%��hQ��	��EƋL�.���`%���8J�)����p�2v�O�6����{o6ӊ��Y��Y�t|QKP�����!q�V�̃>���̠���߯�i�P�W�͚��؛8�h�����:<���w\�y��Ri%K�fQ��T�ʻ�k��j��r骖�'��@��N���TuC9gλ)U��xb@F�0c2����Q��T'F6���6�τ��ئx�߮u�+e�kQx�#qe!��?��]s�-� �6�E�Z;w�p���u3����i�P �]Zy��"��q�οxGs��-ŲQ�]v���λ�����/Q3�K�E���'ɸ�*Y�N̡�̹W���j�y�
p�@�ll3���;�0]��5tNo�o9�m�Hڷ�o�, �9��nV	c�-s3���:r�w���ԧ�=#���Y�JuB3<��$��U6��Q�4�4֧v1�v�X�&_�!KQ��Dx�9��%��i/3����AH8�ZW����;���(Ss�e���47�m5�u���`��-	��f���u����-w�3'x��Y��L<h|���Cܪ�����Ǟ��Z&��L�%?�_�"����p���}JBG��#��,+Lk�� ?��~shvq;��Z�&�
%Z���_2OICp�
�!�\��I�IS|�YU���f����f��5�{�TM#�ʹ<��A�1c7�F�x��)��(���Tʶ"m��~�`�a�J`(�o��yD!���V	r�XI%ӤK*k8z�s�n�3y;l���3�<�xϟc���C_6�ŧ5B�mU��a;��`�-a�OcR��u�� �8lpQ���DU��� �|~a�l����k���Wi�����:�����5�[�M��C����a�>�V3�j�����"D_�A�������h=-���2H�2��xD�,�"���	�D �Ń�hK� �*\�n���x�3Pg偀,@�Zo�h4B?��l�<���m�N�b�E�TY�ٞ{<��p�+N��/;���F���9O-=]�A����^�4"�]4o�S`�,b
�
��;Dk<��L/�rfnw��DrW#5]�D�h�Q4�"�Z�*P��R�����V�� U��\�-��V�B8g�F���}��Z���4f�5�%@ ���o��0���\3�X�xjX}*���*�p�Ih�Njĝ#qxU](�����C�(�>������T�)(�t�M�Ĳ,�ur��a�����p[�`�Z��s��epѼ��1���&�ҙ�!F�46h�z��a���pd�Y^��5c�ZU�ӛ1ʟ�񯉉χ$�%��0�y�����2�՚�=��hp��WR�d͘O}�e~�}$��]wS�B)���s�Ԡ�B�a��it�hc5�p�(�&J�z�X`h�#�J^�9C�MP��Ct��ާ�.|�U\��Ḿ@�N��,F���!j���/�2�5�ɓ���j��-hd���籓*K&1�~b�=�T@켕��`��";�RP��K[`�CbXB�(/VzT����hd>�O���qP�ߘ�Ș�� Ј�K3��!:��[d��֟4	G���n%�����o���KpP zk����e�3≉Tt���A�פr)�חE�ـ���:{f�\�}m�U�v�(�y�ݗ��˒��L����M�iij����1�7� M�p;�~o�ص�9�؍+SB�����K={U��,o5�#@����濲=\ǒJ�Yq�I�v���ZM����o5��� ����X�7[�2إm7kujĘX���n�l���h�y�����H_D���(��_ZRp����OB��^
��E��p˜��x��aԗO`�멂�{��4!���n�H��͗�k���z�����Ro6;�q�P?ш�� MF��6*�������[*į^|[xj��w�ybnH.Cy �.�3ې�u� ���Si��a%_�ѯ��x* q��.�k�U����y��-y�`!������6Zl�9]�����/�	=�qu�b�)�����,��@���#;V�i�Ig��a�h��x�gų搧��p��4�v�m/#! ��9���i��Kvp_rJ�~;���įJ�$�)�͹�:�TE��������3���3�uH4���������,o�Aȯ�1���1����z���V���J���1�Ǉ��
�Q�:7�fw�ǡ@�������Z���a��$����*>�϶�Ul�=�59!²��_@�uo�m��zi+�yO.�n���(�p�y��� _�m��*���1���.�yV���a_�����O�fy��zV�<�Z2FWt^8���U�)1_=�,a�Z�$�iPC��j+��1$G%�F�k�ͧv`%�n�M���<<%N@!r]񆩰60f�����~�ˋ7XlxVHYEB    fa00     3f0 ,��-��;^�⍧#�qqH(�OnUD:��Ol}�֩��:�D�#X��������F�_U��\��
6������;���{v���$��Q^�"�Y�S�W�7��y-L�v��|�Ё;X�n�-%�n�Q��(��
,�As�G��%̅�mWȩ'��c�Žr5Y�����x���z���AP.�1|!�'�w��R��کeIx��o{��m����d}����$�����0 sh�
����Ҿx;`dA�ݖ5jHB��;ܞ|:-{�
��|5��Y�DY�a}(O�XL �S�!Ŗ�ލ��c�h9}�ꈆ�R�s	1`��^�=��J3$:]7��Gh�q�,k��d홆G��N�U��({8C
n����v���Ĺ7�
�?��{"��a��,�lb��|r��,M�b�\�������|ܙ}f�>ՄF-�z4j鬂����i숳�2�S�.E���.p�7	��Uؠ�5Nٮ8RɆ<'?r�o#�ֻQ�Nޒ.	w�x ��;�h�%O�.<�u&�`�*JC�E|Ky ymY��Vr@�y`���f+X��>�%�ʚ`�oD�n0�O2^�	.�q���jƑ{~�xH�5�_(�m31�Ci�1�	��V��j��D]=��aH��̍�����	}�t��i�1���L2�S6�[�t�u�T~�JM��o�U��Xmԇ����)&Q=���ަܢi���2Q�i��s��D���vgNѩM�1&f1ypؙ�9�rV�O���Bq}53�ƻ⟠8&����+u��5�9W��Z7���;��?�y~{����$���T�lP_���,S�1@�ڄƑ�j������ �w��'�X�`W �j<���&�2'W@��b.��x��}���}��m�)g����T<�n{�2�]�����P(+�,�/�s���dwT�H�7LT��W"�:j�Wc����H�;�E6�*��J/­]J�ә���-w��u&DL#�S�����v��:XlxVHYEB    8096     b20֕W��y�R�=a� �[xcz�g����a'qc�*�����d���)8T��ҡ
�O��m��@��"+�OV�G���)�Mq���p�9��*;Դ?���2�jt7~S,���1����s��1��\�x�,��@�r~���B�.'�@7���X~+�x���͡��*���>�f�[T���ڏd֪����g�T:R��9��={�rQxW@���{�/8H$b��?\�!�I�¿GKRQIi����I��eo�Z,NX2̞h��{�������F��e[#v�.Ɨ�?!��E�R�!�+����(���=z��P8��x�X���`(���n�i,�o�p;�?��hud�z��zK��������_h5� ���ؤ���'B%7��b�AV�F���)�Y���忣�4H���#-r���rS�e�Bj�Ik�+�l�܋��[�aXa�j|�r��W5ʮ�֖y� ˜������Y8� ~e1����HuC��"�d<D(�g�i����^�}F)��ī�V#-�oi�RĤo��D���+�J�V�ʹz��������)�FC�ﮆW+����j� �Ã�`f�D�����o�8>�hj��K@<�%l��4�3�����K55*������AH(v%�7y�1eF-���g�.�G�r1{���c��o
(;ig�`����U�W<�KC�g_ 2�=X��z��%��nܸ`�d����ӚzG�BU��OY`㇘䪡2��&zq���b�þ�8����+��j��v޳t����T����㶊��V�[��bE�1E���'�Ҩۯ���#&�l����> �g	�P�x=�|�[�˭�._=}F�F�с�)Â�;*�N���2YE���yV��ˠd��w�� �ډ��II{ױ_'֍�d	��W�!��0N�`Zo��0�؀e���-�u����P���h�ɌOr��݄BN�ȣb
}]61��A��q��&̜�	�	�4�q-/9Zc~Ս���N���h�4�n�^��R���y�qJ���A���l�_�9Vյ��F+�Ȁno�Eؼ �����Ƅ��lY�H�����&�/[f��^����%���J��;��!.�@�HF�R��[�u�96|��P3m+AT��YQmL�-�o@�s�G.�?���?�80�#�5�o�e���tڌ��Ǒ����w�c8b4Dc��_aUˍ��q�R��85/&<G,��IFv�>���X�@�\�b��!8���Rbz&�hv�d�=8{�Vw�(��_��iz�!%5
(�q�P��m�K�s${�ԅUӽDlI�zm�`�b�$���U�w[����s�yta�T��m�}W��Q��ypwJ��Ux�U���3����>�"�+���z�Ѫ���7��@�����Ӕ�u��6��n������ �K2��Z�l�q�֫;y  n���r=<4+?^g��0R_��Ky>��ފ�����z��E�7;�e��ˮ{��Զ�Qy�C��+X59}9
o�5%����%f��$(ds�jy�3��L���N
}=�r�Cj���3V��؎A"gG���O��׬�,�ď��Ÿ�'Aŷr9
b˩J먧���h�Q:��V���N�tB��M�����C0J}�[������lS�Z�`Z�9��N�1�:#�_�4
��	����ئ0���Q֟�!564L6�:�[�z�mR�� </�l3qH%��6'�|c��� �ą¹=;.I�T�+B�����.���uB@����}���q �7^�L6�Z+p�b�����O����M�t/Ԅ6G���48��ez@��9K��Y�[Ȑ�V�7�0���R����h(I*�C)����c�Rz���ۘ��dЉ>��2���g������\�QuLO�Q�\5��� �sp.�B��{8�u	G%�����'�x�m&)]�4�D;�l�����6����i����d���lj빓� ��ɕl�m��v��b���wC�F�័�a�ۦU]LK�9���S��͌9[�,S� L��(ҏ")9��ﱳ�v��U�u���ӯ�w���e�sq�z.��DҪ�Dn���v�����^��{�G���7�y]����XGsP��8��f�On�V�LQ��2����	�ݦ�
17�A$Yu�af�˪�Xڀ�g%q�
�Q�m��'9/w|�.�7�պ�o�Y���`lD���]�����'(z;�ȍ���͇S`� in���h�z�l�c�t��T��z�ɚ:i�.[A٥ᤶ�Jy����,�M�y�IG�A��lA.��.C�B�`:���>:I|��\��Yp�M���?_��؁M� �)���Q�L<�6a	��ݗ�$�=�/�
*_K��ƅ�P��a�f�?����3�1���^e��.���w�6ʥt�(���q��C,;,�!-�ުI��SDen��㫘�aW#� n�ܹa�l��)J!��>�qѱȹXa���5.K^��+��b%q��%�6����4r���EX���XO��PZh��j�X6,���pW�����������`U{PpSR��z�ωb-��I�>����#�d�~-6# )K�gQ��6��)W�s�|M�B{���~;��~5Y��V,��C��ğ����(�5��z1�νæ�ӏ\\�����K��U��5ɽ����.rk����
��qK�4�,m�s�Yu}t(��l�5<���v����8`�DOr�s�	��0"�>�< o3�����3�_x���&#HB[�T���Khb�ד�\�<N![�e�