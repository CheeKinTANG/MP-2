XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���׻~F�)��N��N�.�i����E����ﳛS�MN���{����*�ȃ�{G�tg���"NԪV���$ ��-\?`�i�-����l�F����s�t;�[H��ݭ�}�ƣMʓ.ve�£���(�r���T�n�-�`f��4�R���F�ݞv�K*�J�7�� i[�`(�(]���/����h��2���t�O��'瘫��D5������<�l��ۼ+�"J���U]��X�y�<
}�PYn�(R�J(*A/����j;pR�L!ހ��ԺZ��~m������O�\�kf�*�����񁾫Ċ=�(VG���
#��jW�n[�i{�Mt�#�O	ys�hф�4�a`,���O��J�[>{?�/���?MO�����c �^��E��&zQ4lF^���v�v�[3��O����g�-Ͽ�w��R�c1�Uyh���U�X����uy �����y|h��/��=�̷&���8�q�z�CN6�f�5��4�)]�Oޡ��]?�� f�v�1��.^� E&��RTC�	.��[=J�32# h�J�ݎ
f��ǐ4S��ו�����t��C����N��+��L���vS�E{Z�f�EL��A_%D}�\���Y����3d���A�r[�]
�3]�)^5v�M������h���T�8��{P~<@ۨ?E�0�BoDq(�`��1��s+�{�~�A(�֢��?�XEn�}gqV��k�[z6�Cb����XlxVHYEB    1853     810���}�bf�4]��;�00qk�R(3
עwYLY9��B���(J���0C�c�A���Ӄ�c¢Rt�F��U�����W�h���[��j��+��84-	Sc��i�e����>� ��!.�$��T�U�j�3NB
��M��{��O�Y�Da+Ҹ��ᵆ�з��wgq9�ޚ�$�V�)�O�3}z=g2E�@�MT������&���p�J��|�K���`!	�+�9�\�뗻�X���k6�<w�51�G�΂9������au�aA��z����:�� ګ��-i���K��r�#�D:~7�5MC�����aр���9� kk��莕�R=F�?	��Y�{������Yd��t�w�VZj|~�����L�������G6[�V��:E��i�A�����ɧ���l3���>�BR=:��ڎ�f��%�I�� �P4ۻ+��G��Z��<�g�߀�Ա�$�lغK�BY�r��ln�޿�ПU��PDY)�tJ����<,��D�ȱ#��8�҂������s|.��*B�q�-��s����eJݗ�ɦb��3�/�#�2�jR�����G�#�ݬò� �?~@�D������������*��H!��B�*��^x���e�'�9W��a�.������0p��%̸z����-���y&FJ�Gy�������̈�U��zR��/ {3̓�O��1Z��vm�5��h�p���:��!��U,8�p#�0F�W��E��g*m��+����U�\�S(G50�N+kY��&�����H�T#� �%h������0�_��s���']N��)DC��@����Y��v>U���@
51�^�)��􌰡q_�u_�V�?��H:1�ц��,������ac��P��P�l�-�V@�p4`m�S&?��
�\_ߋ���e��~�`2��8��"�B��*}��d���6B�=��t��D'9L<`�K�g��!)�H�՗g�yA�%�_4<�`++�x6�PtP%3M�`IT�jɫ�Wky2����7>��\�"k��^����|���)+g�k 枳DVJ�06J���8�m;A��w��z_�B�(N��Y����<ӹ�$���@��R��.>{��%�Ƚ��JKGO |B�',��NEo
�!�ζa�5�.����@�Ⱦ����>ӆ�E`����"W��5����·�g��ɮ{K>�e��3H����'�eݍ�K�#-�?b�]8�È6l�D�݌�6챋5y1�!��4@}����ќ�4G'�A�A�~�sJ�xvA��K�~-r�@&�1'6C�%iY=�v)̳R=]T|m�ʣ�{h���'n�,x��X�cCE�)..���uo��)��P�:@F�W�Ar���n�����y���,��u�&�֎�'�6��=d�a�$P��%n�ׯτ%W�(�hAe�����%�l�7�I�/'�c5��g$���f�
a��|Rj����s�j�SK�#�m6?Dm3�n����<>m_&�������Ou3�,6n���q�������&���Q���%�*�$�wS唫�La�00���z�-��#,<�Q L ��WS|Ǯ�'$e�U}gf�z��_�֦�bWYS�޶¾�w��!��ֈ|aÐ�z��p@(%%R���a,A��K��*
0�0ݓM��Aгf����|�׷�x����:���P!�Y��v������6׈�\�F�~��UԖ�����y��&�Xb8'���H�3\؃&�L[F�В���9�������1���������6��Vv�w\��;4|���A��W͘���'|73�{z�"�D-R((V��+l�Y ��d��_2�j���y���B/�^m)�n�;3��i��_tMq�_Y48)�cE�'�?A.����g��U�Q�j��a�gLr4��<��dge8�Me��ݵ�+��g�?��U=`b��,OGb�T��4�r~���Nm�-U������T���M�Ǣ�3�
����g_,��/�n�N�����8�Vԙ<#UJ