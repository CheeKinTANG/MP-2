XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����°'(N>EB�8�}[�W���T4ɨNJ\(atPJ�Zh��R��d�<+���T��@��s�7�^�ੴV<c]}���D)��z:��V������i3�H�g8��l�~r�"�����vc ���@���u�8P\�7�J�_����ʒ��4�˻�'��J��9�BI��JE,ؓ��{侹�?�����i����I�|0���2���dԹ��Ӭ�� �e��bl�e�nA�WNP��m[�����Siciv.d�3���Ȕ-](_�񲖝&5%��d�&�Y2��W���������aU��Am,f�e=B��������P� r��$�=ܧ�r8����ԑ��7KK [���pqô̇�A���>��X���5΀����f0< g)�6G�FДOǾ
�Il$z{��T!�'�c4q+CjE�U��r�r2�aR)��8h#E%�h�`P�� ̀�<~ioG���S�#&@ԃ�d�%�Ϫv�h����ɒ���^��*nd[%��J�O̎�1ȑE�lvNv�#�T�t-)$Ӣe�;q��L�����q6��<-���/�j7���j�y�V%[��s�e{��D�3��o���S*�(�F�W�b������.j��m�x��{�8M;�}5��T�rZ8jp��Չ���)ڢ	4�W�sA����pl�����������RI���$0頋v^�
�����&���=]2�>]5�3Z8!2�#���
	�5��ܭ.�=�z�J|w���ҫ0���XlxVHYEB    6315    1790JF�I>WIgu�`�472��n��
2Y�UW ����}C7���μx��j*uo�A�<{K+B�IV.:P���xG�c�2�a� �R>�)�c�N	���v��vN,��W�%�,
w(\��\�l�
�~�E� )�R�b���H,�9/�������\P�7��?hc=���P�G�dAAO�g���1��y�uI
��?��V���P�Ɠ��W�["1�T����gL�m�����*�:<��2SZ\�������e;IQc�wY����Iu��y�C��#�G#b�� "�P�ef�l�[���{7�B�Ud�l�@���)��nU�F`~��8)�@Ra<Q�g��z�>�]�T^��z��	{ZV�Y��8=�(��,e��r�B���`���<�e"f�g7�_�z�myP~8�X���ɳ��9AEw�+�\��t�q-5���<��O Ո����vRhr6=臦U���Y�#��8�c,\8����űF�����G���f�<u�x��DU�!E`��<��[.Ew�N����1���y��_Q�ss��z���b�1f8!*;�����<P0y!j}�� 4�f�pŪ\�U6�p�ĩ~dŦh��3]a��H1}��,�G�ߗ~7@�@�z����r4`�RlG�wCcy�|p�قós}G#�����It8��]���*�H�?�)���71Ž^���VH�ܟ�(� �\&'�HX�#>�Ux�[��iFSʶ��$2���I55vf_̡66�K�Y|-nE��G9az552���| u���cgHG\[�e��g��Q�[�b�߯����K<����T=�&n����%сj�[�<S8�o��n`��O`
��"UJ8���y�0d/)hN���,�ohg���p��Ь*�V������p3�E��Ԑ���2�陼���T�.e��"y�G��k�y"\
I7-ŭ���5 $YÌR�?t�hBˠ:�l1���8ivuCH8�������m>�T�sq�j/$���0���3�`;	~ � &�-#�y��r���?xʪjz�����?���{��!25�,5���W ;���ZT�hYe��+�"�>m�������z�HǬP[����������*����r�.����B� ?��V���=�B���0�:����_�Q$�ymR�R.���Ť���R���1+q�ʄ��{u7ڑİ��ޜ1`:@��mJ���72����iboJخ�|�j#�6�Ri
7w�I�7N�� ������<HT�����u�G`��߷^�z�$5�A����X'���4@���PkN��@`�U�����n�9�İ�]�x��d�sI_��Uܴ-9�4, ����n����#��i:�)�D�We�7�Q�iz<c����*�&%K�)�x3nʭxNRn!���k�$��xs�3��[�2��k�	��o���R����:����	���:� &F!@o�q=���V�&;����L?�x�b�D�Z`�Xd�Ky�YZ);�B�@��R�f�Ԓʸ'M#�M4������[չh�����X�����/�-��O�C0���$�=������k�S�q��=L��@o� NY��Uc����n��ND��
D��t�æ�D�U3�o"i;S�W�ݿ��`�t���$ǌ':_k�/F�?�5�P���~��%����Ҩ�~aJs[��@�C��G{ ��zq��ng��?��YiE�YA]�k�>����ə�<d�4;&6��	��L� �E�%�G4��@�=a㝦���1lk�ȸ26[Q��jd�C�Щ��IA$Qި�e����Ǒ^���N^(I$�kd�?x��e���F�?(�xX3@���oL�f _7E)Gb�0�A�77);�W`�ab����mv'~y�9(�[X�=m�G����`���f���q"�Aѽ��<-�B�8�q�XL��KG�w,�8�#=x#�%���:�NZ�p����%���1����B&~�nm���P5>3�K��*;�e��9:�۟=� L��X%v/��$e$)]{���E㇓�S�|)���$��+�3x��vN�.���w��@�F�o���C�qZP�DvՁE��*�M�4���Psj�3["@�0q ��ٰ��Q`
�l��x1����`�1�gj�$��G�� �CR������l"4��4/5ґ�J�h�G�Ը�iK�%�IZ��Z�<�U�y^�����s�~V�32��|��e3�
�yn�
����#�_@�?5��7�9��'VI��{L-v�ێ�^U`-|Hq2���O��a�E~��uB�hh�^A0jd���+/��-k�HW�~��k��*�{�2��mx����h�Bֱe{�U5�h��r�k>�ya7۩*JR@şZZ���o�E����JZH
H��L%ng
����ʔ1;��nT�4��撨)��F#qlN�d*�|�<e��� kѢJD;�&�f�4p��ٴ���� u�tu����CHMք�v,��jA�'J��Ѻ��@$ѝ���꾔�>^�6ht��vh'���*� �u�M\��j��������v�9�Z�1��Q[!^5���U������ou������S���8#X��*E���:r�4��3����E�p>.��m�b�0��=�WBU�cA(��yoe�3�����0���
�T���(��
��p|��;WȮ�=�TR�C�b���� �=����O8�l�`����(�i����T�o��Y�ʹ�mG��N6��c-NPΉ�i�״�)m���+�^���@���]��ak�#.Q�CB\ޯ�R� w�����OZ�l% �x�g�~��D
c^9c��i����9�Y�����I^����� ��~�$Y�I�-2�J<��q+�P��:8��W��`�8�-��U}�'�0d��+)(�/��%U�u�;�ca�xF2�k%��GSc ٙ�|����R��h����s�9=v�$h��X�����iH��$A��D���N��1X�H��=��ϒA��d�� ܺ��n;��n��OM�Ha���8��� ]?I��������ѐĕ���n=�m�٫׶�-���:���3w�)9=F�つy)��-��D���[���%�>�n���b["x✟��,^�L�
tf1*�ɛ���F���?��&-���׏����J�s1Ui~��b{2D^z���7\�������uU��)�����Qa����)���H�􃠋�/�z�lE��6�{��"�m�A����Pw��a�rZ�A�ߑ;W���r��m�}?f,w+�
�'Z�!	����
hB�x/�����'�\N.���.��[�����?FM4R�1T?�z�#ؗ��2u��+wg5,��¤ڎu[[�*?j.�_!a��s�����rV:��� �3'�ϒ܈����Vʀ��r3M^#�;'?����b�v�P�9����<�砳_r�Ҋ��tL���e,X���=6<9ɒ�ѥ^"{�.�ɎH�t#Eum�!�F��i��YO�W`�4���Z8M�:�H��B��~�fÊ ���
�ȱ�[�q.�Ş9׹A���V�y�-zp�ͳJ�����x�|�~�Jwn9��K�ț!�E�y9|MsŚԎ��ӌ�X�1��C��C6�[�ooS��#㗵�蓶5�F��$�̓г�zEK��1m;����џOra����c���N��b���K��ǫ� T��o��v�����Y4�M�Ǐ���;t��p������M`ugh�W.H�|�2��g���l�
�X���7���\�V�(߬cR	?�@m�!�� ئD8��~IYT�*FԽ��>�l�����wR�����(��o�s�����vωNס�M�=��#��?���3�p��|�}�wP����2+��z����+�E`�Zq ���β�?sVA��m2�$�D�#D��ֶ����YR�a��Zh��ti��x�Q9o?����\q�o���Vx��I�}ۡ�fQ��0:>�ټ�%�stܸ�%X3i�&F]�4�]�α����a1��kͨtC .iO��ky�8���m!o[;R�'�5��������?%�}��G�kM�&����������$$^;��-l�<��o��BzN'!.�aN����T��7𔘸Y- �@Z('���ax�QqG�drN��d��A �wL��4��ۂb%�ځ�vw�>x��>!�'�����}>��,��,*�ۮ�k>î¬�6�u>�KS�R	� *U��x��q�Uv��c�~;�2�Zm�0��-֠%�#�k`nY
�)����e~�|��r꽙�?�E}�6)��1�/Gw7B�
{�s��L�zN���8>�kb��_ն`�aZ�!-�R�_��A7:�@.Kd23Y�vq�����'��Ԭ|��ؓZ\�,4o����GdX����{X�#�t:��X(�3��.��y�S��B��o�3���8���'� 1���溾�wƐ���ݪ�����=8�����݋��+�Ty�RIܯ�`6Q����(�Y)��y�`/pb�V�,��@4�s�;%���<-��F���2�z�R�No���~������y [ې�����N�f�)8�'H��C�n�E���,��%sdx������E%/��A�
#fB�rRN��Hʺ5�މ�`�Ѣh��{�ܵ`���cL�ܞ��~�N�ַW����ܒ�9����E
qJ^�|����h'<�㥦fV���fuP��e�_�T���2C��	�6� ���^&wЊ���N�k��Ǳ��w�" 5(����L*T��Gx�e �s@�����ό�r�!�4ሽ1y�A��LD�;L]x�>�zp
�"�:g��ɋ�,����V� B�._��E�q�i�5� (�����Υm�Ԩk�RT`����P��:�v2�XE��vȄ����s�O��F��U��:�����	�H9��;;6��a6�ܳ7$��"������|�,vRLvְk�T]��hg�Bc�F�10MA.Ivp�-'��L̡b$c(��3E`�(�L�b���Q����@90{�&�& #��jg�3��9��y)&d�U�T�H�>�,Y�d-(꺤�5Zk�uk����g��h�І�qB����� �y��%Dو#�|*,�=�,ӂ�{������8��s�L�eE �oa�V4�!��YJv|+�pKbr(�#�x����I�f}� k"8
�2��`}�_��vH����v�r��>dCE��U6�I�H�^=g�Z�>���^��gsmx�j5Bԁ��ֻ��{��:?`����O�Ĭ��
�0a�{)��#N��춁Vh��^=����MS�����$�����Gl�F4�I�>໗4�o �֠4cv��ǜ� �+X�]jՎ�SP�E�Y��7��q�������~KD[�cvm%ho�Q$�����^�R[�JP�k@��Q����׬)�x[sц�8���v*������`��s�B�-��i���T�N�J�<M��K�F��Ar=��C�W3(޶?.�Ejͭ�y��bn=�oێ.{��9���Fo��7;�yAv�mΈe��oL&E0�Rt���lu�2�.WU�LYPJ-�3!��<�Ӄ�@u���9�N��͌�@�'�l�t�{ D���쾺���KjOEh�(�O��*&u��ӛKy@�{mn�}{��Έ*�EB���/��""��!*�ବ�'�n����02�L�I	�n����HY�N�Ơ%Qsf�i-��o'H��<��<�l�|����yZt�#����KK�s�@]�^�u9�,�8��!��of�/O���э�tAt8���JED�C�K��o�K,��G	���QM�����Ƒ���F�7S;2n��G�T��Q��p�9�IFhJB�!�$��u! 1M��qi�s0�CbG���p�!�;<Lv�r�`DH5z�x