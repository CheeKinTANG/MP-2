XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.�"�c�N&;d:A �\CtOђ6��.���J�W%M� �O�
��pچ��}j�ΰ/�cR�
��k����_�:O��9��&02����	�s;кy]9�p�R�����.���5�F�i�'��ZRR�/��1�w�C����4�?}xv~e�X����m)84Q���_����i����V9�S�)���9Vi}��-i�"G��|��,��A��ۘ�м���?��� .x�t�P��o�>���z��|�ٳ\�2�&8y����@6�Hm���	��y���a�I ��Z�m	��gP��P�<�2�=�ҙ]�c���{���+�k�����,D8����us�3�d�Kr�5yk�T��0�Ȱ�"�q����$��R>x���)P�Pu�Uַ���đ�!ѝ$���c�v.c��,d�͘U�K�JB-���x=՚%��y��驒c��#Z��2��k��;�T���]1�Em�B	��È7c��ӥq՘��_��eDЦ:��ß�V1Nw��Je�zq�kV��Y�~��e75��>��
8�4�����v���4	��K�oT/>�I�v��Fh,i����Cc%�æoFGjoo�x깢UQ�^������ߒ��"�!TWmD�Lz?����A�̙�ǎ�EW���6�5I�����#�,*.Q+���	�cL�FD�7���&���26D^W���ͦ_�
:z���&��(��Q7���V�2z�S,�/m��.�q�eXlxVHYEB    1853     810*}�;��թ'���`�x�ᵀ8�x-��\SV����:���p�M!GJD=e�6��Q���Ex�P�_����y��Yf)^���̵��;���xy��#�	iQ����]XO�<W��YȚ֖�-$K3�j�y�#b!i*;R��ꬳ�Y|�BXnHm4�M�5 �jCD��/#~܎�+/�TXz����W�boٗ t��Ί'�SeF����A���DsVh�c�KК�:�Y����=+��'���+�{T�`I=����t!�R��0Z�r�T��l��Nz�A��`.���Z�q��!'m�7���_�3Dr.�{;�v���u��q�����)>�P�� �Y�ֶYQ��+�s�V�I�à(L5{���"���!�,����gqGNVw��:x����в�/VB|a�/#zY'� z�ڎ.莓N3$���J����]�'
zSOQٓ?�n؂s��N�r�L��BC-��2r�vr�5p�d���؉/��R�v^h�<���wb3�0���4.�A�ĵꉃ+��1q����N��0>� "g4��U����.`���%�èХ�7��O���JZ���[O^�>T�M��;:���0�Y3
���\��R�Av���f��8�d�T��z0R��;34va��������F�5d������P���/՛]�ѓժG��A��CB�͛C�e�WHU����:Ft+8��zU/{�,_�ʴ���N��b��m���6���d]>�"��e�K�d��s�O�!����6���3p���*�1��@�6� Y��ad"
y[�UZ����T��3�sbH�m���H�����'��y3�k�ǫ<����9J��Kgk֠W��(ȧ��m1�	�i��dh��n�itRj����I�p�W�q�����`G\Dc�aD_8���5fI���mE�j���a��@+�MMRH�Y�(	r:���k��C�F�]=�6ܣ������&��1�1of�\��a5� ��c�,�*���e�D	,�O��1�%�X�6�ڀ��DF+H������b ���OFR@��fl�Aj�A4�T�w�=�}m�ko�� ��.�_��^�����T�6���H��x���ȸ��3�2�)�SJ�����q�,6N��kK�sBA��iW	�$��N�ݞ:�����;��5_�Pˉ��F��wF�up�� 0���n�;�ל���5-gU/�O�#Ջn�Lћ�l���rAV�� Dq�݇6ww,u�С@�D>}�L��]7�İ����[�[�y�}6Wd(���(�kn���3f?�}��Ҵ+~(m9zB P4w���<V,�����!2ȔQ��
0橆��D��s�z:�1��5�����x�9�W�°��~c��j��2��[2ޟ�B9������ۆoE/��B�z�
�4S�m��H�S�*��B��Ĝ�����}5Q�p�M|�U�Z���U{Bg�"9#���MD�}r�� �DN�C���#!}��Rv�*Z�i`���¹��"k�$�L�HF�k��=<p=�`��`�n�]"N3�QK��Pc�ޚT��v{�껬��?߻zV���Ns&J��A��:,l����{��l�2_z���B�i��{�~2�p�_��	n�1���OmǇK��Kcoi=V�+�Y�W�+��|Ŝ��R�����0Db��Ar-��U
��:�l\Bţoi:5>/Q6��e	v�QӉ=��E����/���4���8CWs�i�;��,�.ufi��w�hꬃ�D�tO(R��M\W\k^�>��c��a[��5ף�=�ke�K����o��> �12؀s��g+����il���8ʃi%�����P'#�zݜK���7+H� �UT|����'�V�Zym-U�h�����!��5���B�͜�<0¶{���$�i�26|^69��e(X��,3m9e�����-��KzJwu5�y泮`�e"vx�J�Ht��d�0��6��>p�S}���L����M�_q��	�ٮdy������?7W�����"��z��