XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o�����D�?�
�F.
��kt�%'���}�����Vu]A����/vl�RUh���e�)���}MZ~q�70�5x-yt�xӤq'��I�5:�<���d�>H|��LV��*H�Nr�������I��g�c�I�Rg�֋�W�R}���	l+������ڀW��9��<	�F2X�dc*4�"~˩�?�SV��Ќ��t��4�-!���\$��y멾�6?M�Oa;L6QRe��W��X8��׵��V����T�*���?am�RY�X��!�w4��9]��^@�w�b�Q^��*�۝<�p5HR�h���N��ۀ]�M�3a��5n��c���A7���>�-i�7���Wr~]�`L}]���jC��i5�T���i��L7m��U�.��T��Hݏ"�Y�fƌ��=a���F-����c��0�\�::7cl��+
ou���δ���S>��>h:T�;,:b���U�wZ#�y�5�сv���5�Ō�RL�y:<ʴ1���ɉy�4���3��-�1������7�$$.�١~�e^�[OE�֙Q+4s'�{>�W��/��\���;U�t��-{����`��hfD�����ܹPE�1[���䟳�" ��w�Dp�m��0�o��t�m�	��w�묖XG���}�Rh�w�Nw/!yL�o@��`U	e����}�v�����a��8�Y���5���7#`��Xv~��B�$Z�c��-ʱ!�F���b޼f�|�XlxVHYEB    da59    2e30@�>�g���&�q �3v�o����2��_[��S��_{Щ
�]b͇�ghM�j��l�c���u�CU���.�_�+�vO@>f�;����ZE�<�A#)�m�Yrn� ��@M׏�c��Ƕ}����)��;���p��Pƴ�l,���u;�\�����eg���Z+�N}��YN�8���\ ��4��$�sL�yGH]�����\`���1�.���f���֎k,vL��ӝ-uˋp{���5���w\�X�V&�u�����$Qg�Eŭ�:_q�q���`�C�Zw��'�k#�9<s�<��S���mB��%��b�?L]�2�M�{p�`�?��
<�{ Z�WfR�Q�ؔ�*�.B�Ko�a�J:g��ײ���R��}�VZ�^�d�2��o�����C���r�H.�*Q�$B�
���}t�,6@��8�z����I��wUz\`x '��i�q�E�5��#Ԍ�������J�܇X�A,s��h�U�Ƴ�mW7��� �Sz	!�ů� {��Ɏ��B�>-���-R�0*�߹�Z��'����<�幑�q'��+h����>�#�m���C��&m(�
�'���{5���4n��n�Z�{��,����ݸ�ڤ�S���xt�{��j�{�t���$�9�|�aX�>��`�{�7�m�Ʃ���u,�ꨲa^��׻O]Xꆿy[�):��mۏ���ۨ7}��r~֜���D�D�����7=�׽)�=��U�Y�"�wPn�Y��?����\�g=�{����P_��/�|w0��g�⎘5~���U6~R@���*��k�Xh��TS|�܀�X����R�)���|-��CS�"�I�����f��_���0?��t&jI	�l^�*k^]h��Iv��������,+E*Z�C�%�͉ &�:�Ŀ��вʞ�ӎv��J-��-A�*�υ��kL3�cp�0ye�ؠ���!F�oGr�������P���!���f4�J���=l	���(Z�J>�v�dH9�&����f�i�!0rJ��.��oX�
D��4��	��#��t�T���F}+�J� Gm�N��B���JW?������lE*�Qb;J z�\��{�����r�ڑ�(?�k�o�I[�c�:�x�]�k��"Wxʪ����*�Q�T�i5����4�h���)M#6<����ro��|������q!>l���͈@w� �c�P�F���`��fW���h�Z#�1�9�}u�C���|J��#�E��ݾˮ��B:��q�)Z�tJ��!d�':����~'��5=9*��KXx��qEi?�����BʺzCE?lR�I�6�`�j�j�̀v�%�����6����:DK��s��el�p�ǯ�%�lL�q�!_lyuX�Ad�r���wq�ىd^OR������fj�aᤛ��i��~��`��l��'w��<�/�Z��-��e%�E��i�۶QC�u��TqEX��X������n���H�F��C-.����K.W�ʼ�	�bcH��ӊZ������%֏��J^��}����&�T'z`��X�^��9e��Q6/qv�Ξ�n��3��@/�,Jx�ƃ�,�~� Oa��Ҥ����A�#�Ԣ%P"���f����eH�'�b��n�[�R���gN�G�O�5���`��≇�|2\�	u$���"�
���#���m�L�S�r��ҹ�7fq�����C���gt���s2��N�*��y4�jȹ�&X4v�1������Qxs��)� �f;ZS������=u!�0��)@��ϵ;������LB��a��yߨ�F����R,�Ҭ ��������>'ci[H6���s��ݪM}�����t�&+{���_2ץ�������۞-Ć-Rl���Q�0\5�G������[~9��OAƍa�6I~��� �ͨ�����Ί)jFm1�
��)(�r
�#y�*t�J\QfS���D�����z�����Oa��D�ؐjÂT)�b����v�y������ț��	�?����^�_W�,���:�ԁ��m�(��n���n��M1c��~/L��z?-u���	�V�[��6{�����C��&�p��h����L	�D�2�������?�+�#�rl:�>��;���2�03��_W8ب��U�-����t.�m��&&�8wQ�k4�^hUH�ގ?����8����t&�҂���ֵΞ ���B���~w������^�4luz�S�R�kq��P�op����IaTi�Hq��I)3ɇ�ƅ�,P7B\���πꌇ���4�$���w>�!���e��.?��]�������(<ٛ���B�w�����LbJ�DZ+�ђR%jf{ ��J��p�a�n�)���+!��[��=�:�,�j�eV�[�9�>sP��^�d�g�7���0�A?I�n���\�*B�>_Ȕ�=(��>׮�������jgȗ$JE\]Sc���s�f�LD�X��<lej g��F���>�h_���k�P�O�t�9��b�����7􌡷�1�-&!	� ��8e@{˗R�_��TuҢ�~��@Ր4���H��rX��x)60�m֦U?�E�$)�9��&z���H�}�F�[,n���tYW�&
:"�	2U��>�A.��NY�Eo�N�b'�| �f@�I3@�D�DݯtӚP��v a�v����]PDYwB"NZ�$�Q��a����5;����x�b�&V��Cq�eh�b�I�\,oc��R �iQ
�J��u�k�ȃ`8���� ގd��˺�'�4%jW}�á�ZS�`�@���Z?V�<J���p*&y�1%ŕ��^(Ǚ�C/�ALBE��)����w�W�|��r܋��Y�g�?&܉��z9�(�����R}bb��sO��r��a���� ��}������{��S���־��G�n��ao�2�(��F���-�����l��R��9 ���szC��oܞ�tbu�������;>@l����~�P+�ms3�p�]�.��T�麑A:3���B�{fR�-����E$���bNl�����>��l���΍��q�%z���0�"�I	�QE�[D�8��n#�O��5�P>;Pc>�Qgb����%�V��'�Rb�J�H��s����`��q���� ���W�j�l���zp�{$�/�Ф��>G���`p|��J��d
͢f��-w�*��kl�����!��2�<�5�,�
�zV6h|{TM9� ��SӺ��

]�A�;t�i+�r ā�ȧ��+�\v+�n��0u�I�V'F�#*k~�W��y�3gh�o �w(z,N���Cq�Var��I���+���d��@;TeG�m���2[F}�Z�7���S�c3D�`����#F���p:�Z���Ԗ����~�#
#/:2u�s�`�G\�v�[n�ٽ�2��UD_PvT��[�$��N��Ro
:I8�!j|�!ע�����-̫�&��沄�X�ĺ�aN��JjDL{��F�wt�^�c�j�*a�Ut���Y�1t_^W�a(��Vf��E2I����jX(S�VC"��$���?o+L��ARXt�h݄x��$m6]�����BH�R�Vq�־�K�)���Vʊ2�fK��k�ܟ���h�V�D]���|��.��X[�	3��+1w��8�?���q|V��Q��^�M�����8�7��%Fv��{�雥Q8���(r����be�'o��%Ax̯��o�]��j"��.��":ŠJ����}0�Vz��X�
q3`���*�L���ʼ�)���8�w3,Q=�p~��~�v#B~{�<��Դx��Z�J^ݼ��/upyF-v��Z�#C����8nE}�k��aHN1�f3"?}<:�
�wݲ���hn�Ρ���g5�[����h��Q/���Z��_�<aYǰT2�3 �	�&��b2��Y�z^W%��=_�)�}�D�G{�(��9��;s�Oh�$��~�l�9cyJ@� I�g��D3����7���j;�r��������\[KP3Y�E�⇹PAF�����ji��e9�� ��)�B.笸y���N��ɱ�?��NG(�����
��-w�\���sB���������#����K~y3-q�i���F�v!ғ�K�:j�u�*�:�����+(5�$L�j�k��\ްF�
!ͮå��5jX"[ڤ�EƲ��Iw��Uv65߄{!ʡ*;[E7Z���(�Y�D���J��B�~2��E��������o�R�ٽo���\VZ��]A]�݁��]4t���n5��K#��������Ku�� _@��L^��ֵ�<�����J��0H ���`��`�^�6c1Ӗ;bT�*����7}��j�x}��R�Kػ2�YR ����P��Z]�	.R���{�E���<Á)��7���^�Z^����D���	�
��~f���E'1�N�����6��o�:>����vi��!��.V��h"�C��a��=#C�#(o��I ��t%S����"���k�	[��#W��щ�C�>O�3룆�yh�����rH�K%�w8z�=�=^�p\�vn�WNj�, 6s@���E����j$�%���k�p`j���MӸr�j�&�,G���.!y�ߺIsv��7��Z8v�[��eNI�JP�e80�����H�J[Uˬ���
����Z��N�\�M9%�SSN��D{�� ���p��9DN�F�>I38�V�M��ΓЉ�� 5�ܭ�
:������A[�>\���}��D��`��Q�왺���C��N�R|�������ȁ#Y��h-Z���o�{�̚�O��k�gF�����æ�cpZ<�М_�K Y�&\�Ka�3
WG��d>���0lQ�����=�W�P%�b�;;��j�r>ٙV`��ܐ��u6Ƞ��,�����BVb��2	�E�P
�4���z���,���&>�SU4�d�4�$����/����.N�$�t�9�s�"���� /�̕�8������N�FM6�98jIN$.�n9��7��}�qȱ�h��:ۖ3��D�Mr�TQ�)�.,6i����Y'q��g��T�qA`̗���-W$O��0���3qd����n�\������\t!��![�1�A�����YtN�*ȏ3B�m����^��ȅ!,����{m��c&l����}1L^+D&�(X�xRqa6�h�^$Ո�lu^�>M�#�W?���7��j�,��  �L�ֶ�%`_�����ה�g[��='t�&FGꠄy�̈́�Q�5� :u/�T#Ñ'���p"'�a�.�p(�m���� �������,�N�������)��ڄ�h�x��Q�5��uD�X�VN��uȡ3֛��:&ʾ_eXc�t9�Vkn4fh7��.p�5�ѣx��5���p3���Vʈ1TqzD����N��Tv�me�#���}����{���3ŅA��pI�p�=��`�}JBoo�#�O�W����0x��®NE^j��붕� ��u�:�v9�M=�{�*41r��qK6c�M6�a���U��hS0��	�~Z����(�n+�s,�Dٚ�):}��;�h>S�*�%�Zf6��R���O���TA�`��Y��ϙL���+C�9�W1�����xj*&M6��T}\�@�OWd��m�{#>[��e��0�"��B[xq�ۻ�����k���ؤ��r��,V6��t��)=�8g�)/���N����oo:+k��aݯݵd��$�r*�� mo�b$33�kl�j�V���1�#I���|"�����1N������d1�?C�>��6nL����ǡ��6@1��>�´4.^��x�r��������T�l��M}x��Kt�xL��A{���OsI?��h���϶y����]�4����>����gq�#�-fY)��+>=��N;
�6#����#35�O��r���I��;�6M߅-©�K���!����t�ɩ�|�&i� +c���u��8i�ͽY�Ұ�
@�Z
���:��������qtf���:#j�\�O�bn��J�س0���C��zh�
|\o���V�Kۗ��?��x�+i[@0����_Cv ��غ������ �+ۓi0pD�E���W&_�������A'�V|�v�Lo�"���Ս��q%6��m!�v�E��w�A&�T��9c"���VMF�粨���&6P�O��5�6[��L��J9��M�-�0R��3}�H4k�d�M)�w��55���s�� ���5J��?�6bh>��G͠7?�zI>����7	�@-�S�8�A䱑�J���f8�h�>$X��#��N�C� П��4��1gk\
�b�n�^��O�JJ����X�mkd��F�}r߳Q,�%�S-��26�ņ�5�E�6.��?O�M@�t��H���������(���46=�Fbտ��c'*����cLy7K:�b�!�l`-�[<'7��_��VKB�Z&�hq?�kՆ������t�����Kc���]Z�k������ ��x&�"$����k�1�C��Aϣ2���nz�=`rbl�,Ԏ8E=-lr�����K����'M~�{���� N��������J��h;	o5�`��Qs/�k'�Ȏ�/�c�bE0r�#��A��j���bVUVt.+@ ����S��&۱A?1�<#�� ���!�����]��dZ�|v{N���r-V&�?>��
��ǲF dk.h�c���p4d��H���=�0�Z
���#5��ff�P/�b��M�%���s�s͌>���1]�
����2�����&��]��'�`	�:}�F�*������l�8�^"�IY�,�ٸ����.[��n��U�� �ͳ�&�a�G3�YC Qߜ�ν]�����mh_����%ߗ�����:ݔN2��ƿBuu�����0o��Qf�U��bl��o��L	ohq�]R��iW�c�&ɟ�~>1�Iy�|.�Y�����C���%:�kĘFP�x�-���xX�����Z�Ut�v!�m o��2���2w�i,�*�VV�����M�6ū}$�N_���c��.�� �_�U:ܺ��d/��<��'п�Ib�$��y��F��:]�N)��iQ�����Dg;d�)��d�u�j �rB��0���A��N�=E&������
�G"�1z�]2�$`Pw�Ê4_L]E�H+�3a޿ٜ�#:(;c�I�;�������:"d�v��\�/N+�S�ד��Cv��E]d���t�zo)Ნ�wϭf�a�$l�r����[�A����8�A���2�k���}tN鋚(�鹅<� {���%m�X�3��m�ƃq����Q���i�lA̐C�^�W���j�+9��8��=WMb�>��\4t{�*npq�*{�h��9��%���B�B��[��y�?�� `�JC�֭�فrl#�ur�Ǩ�鲉 �q����[�(���&0����I����s��,C��S]�Ǝ�A| M�k�t0'e4=���9��Zo�����u�_l��Gǫ����ZD=�u�����#�a깩�G�G��A�y�ɹ&Щ��h��$���������!-����x���Ң�����\���Xt}zk���"b
	�a �r(v&��+]o���Tp�f�Ї���o�_��/�0mp�
�䯪fmȎ�|��6���rH�1��VuR/�I�8uSDo9{��t�����7F6�������������Q�1GW5X�����}�o@�4{:�c�0VF�����$N'���]���3]94�����>̽*(�ȡ���+T15y��8������H��$���"z�oT��/�-A5z"����'Ǭ��D�!�H��Lo�U��� �K��H8Rs�S�}*�Rд���}ͺa��Y��{��%�]��q�p0����F�ك�~���ݼ�klNL��h�m�[��*��C����F��M%�B2�YHwVv�����d��*��S�xm/;|XE��h�ʭm�h[ʀآ���_��fH@T�Ğ;����aS��E��F����:��|�_,�h����������2{4�y�}8�kZ}]5W�D��s�ϻ�p���UԊ�z�������?Ɯ��<���2�1+
���i��-�&CܿPBI����6Sy���d���N Vd���ښ��{s\�yx�m	H��P�� z�U�F��v�X�m�xoԹ�&��e�띾���J��6,��h�� /L1#fCC��G��rRr�|R1%���:�����襪KlR+=�I*O�.��3�%���-���^C\���N,v��>����)E��-��5���Y1��lR�O.,��RO}@_~���N��Sm�C���	Rv�{QJ[f._1�3CGNi��؂`}`��b8Gb�m4g�3>Y� ����!�q1Ŕ �o����'k]��;�NL��oK.Q�X���~M������3j]�A��d�����t��"�^t^D�+W5YS�g�!������Ms8�� �El�\!��+��ٯdo��:��pP��P��Q�$�7^�G$�li#7Z��|}'��T�t��Y\��Q9.�A�5�@Wriq�p ��Sؓ��B}�O�m�m����M�����V=ޯ�+t�mu	a5��8��e�t�g_��2f���nEN�.|�.^�i��s��[��rI� k�0�������B?��q2��t�j+l�'�8�����K{W�����l��C������(��vg/�a��D�P&~���v���_�����)u+È��ݷB��&p ���{�ڇ�qL��5�>7�_Քj���txP f�Y�k��!N�j>��j�P�T�W�$_ز��r�c;`�~��-���O�U�۴��d+�w������&:ę����{�L{޶$Fe������7��?���H����N.a?���q���j�fV���]Hv�.Q����7?��l��J�/^6� #�O�h������َ�Ac�>� ��1ᡥ��(h�L�ʆ���)�MF>��Vpxl�ݔ�޾��8ݻ���s=�]c�Wr��r�dQ��>p�Z�`��,$�Y2:�ҩ�>���"1'du��2k�mq����k8T��N�~+�h��e��Y5>ϥ!�3����D���+�힛��֖:fIT����68�M��(��2�%s��Y{"q����]=1d���n�Y�W[�xK�m�i�oe�z$N��t�>6��Ds}�\;$���hE�\���f9Ze��U�Os�P���/�@�p1�4#���� �km�������@h�#F���΂����w���*�7㹟N�Ґ�5�9�U���}&r�T�I��_��d��X�$���*�gEn-;�*=/�.QA=N<I#߮?cL�{�&����P� �[�Q�j ��b���5	�	�"&B��c���:���j0�/���i�~g�+���p���Bx��3v�VH�e��a@���"����x���rYW��E8D}��]�ƒAmM ��_+��0�1����6k�(���N�H�1ԹjT[�Wn��vߓ������E$k�fp>\5�{���e .=��ŶYU�dv�z����֦�\�˶'O�#C�+vB��z{݁�'�lJ�G�<��a�3� &�5�W��0�w9��z}��Y�'�(QKs�,-k �m�Y�P�TC-�<����?���=���0��������Hlg
��~������Xt�j���^fS`������B�D{��^��9w<��l���\6�SQ�86`B%�����^}�>�>1o�
�g``s]��`�=���5kυV�vP��2�2�v��*|��`s�&]�I��ﺒ�4k3�#�T������b4t>���^Ry�_Τ~l	�oe$Ob|:����U��̔� �l�މ[A�*�~��&�XA���8T$�5w�EIV���T7��UXOT�3�\�J�Cz�L{e(�C*8��/�4|5�ꅧo�ws4�?^�D�OS�������� [�Trj`�(d�AP@��q(���e�A��.�������q�<g�S��7�e�5M!�"�p�fF�9 ����f�z\3>��F*Qx��h� ��+b'�f�Qo��r�w�CMO��ل�1��w� T��:��H(FP�xS�^G��N�J U��Ʀ������nʰ��'Y����v ���SE��nCv>d��_;e �}d��|,��~�0���R��+s;���Zn�׺�bA��>]�RC��u`�/'dp�z�;�a9F;��<�e!�z+�{? �\�	�s�ٱ]ZJ؈^1;
�U&��ԣ�y>��P����/���#�)�LG厂 ��}`���'�sxHw4�k�=����_o�Xy��YL��j�u;ܺ*u�C�8ގ����&o�	>5=˰4���Mu�v�8sz���Ϥ[�	>F���V�E
��ϴ4���v��,R��fR��v�����h�m�_D�.V���lO*��Tݣ���
��@W}��U�l#q�������b��0���9���5
y�2�N
���>���WCX�}D��T~B&�L���۰
L��D܌k���'I��5��_�d��\�W4�����.���S��y�G�X�ܔO���@[O�����XE��I������Em�[6��@�M�Z�F����~���	�����iH֏��v�x� 1��ucϘ�����7{�m	H�s�O)L[��_k�3�(Q�(|7X��?>�}$�b<	�s�Q4�F(Ǳ)�Sa�����0����깴us
�}f���P�yaE������ehH��V!������eyA ��9� ��k8Z�Ẋ�jy!'�L�9��2�	�{Q��H�����������QG�_+�|*$�4����"
X1['�HE��2���MN���2.¥�a߹AH1���A7f�.��Ą�_5�?���3vA���%�{��~�}�z��xNp����W/�˵
(�b(�Mb��}��%��o�4<W�_��aǛڴC,���N�_����:>�A��~�D�o�e��uXm�K7o��V�%W\!�4:1|!�N؆��Cf�rfh���r�2�I[�H ��,k��xp�W�X�Z����GFp�P��ʋ����g�AT����� Xڰ�E6�I�qv����($��[��5�#[%��G̜�Em�9�ҙJmpM͋@]�mJ�|i�j���?�P���Q�b������wZ���d����|
pF�9����(���(���KSZ���H����_�E��.���w���T��95>Ĝ�M�T�H��R��a�h�FQ�x�����i�ZK�g�Z�N�!�ێ��3�a����̄�:2�����9���>fGT5��h�h�x��{3�٣�U���<���S}���	���$���P���>�-ar��tU��I�x��Og��V�:ψ�;z���ygd��P��(�h�!bW�ᙚP̧��}�R��A�[�Q��ϋ9}B�6{�>́noj��TVbO�a�p|�}�!/Ji�