XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ѷ�� ��1�i�9:	�G����T�F4~ҡ�����bO�ا�g
+E	l+��A?������fE=}��s�SE'���� ��qZ�<��~�X�8�v,�x���sʐz��c�^0�T�D̼2#�Zt�)��πB�N\Kc���#�b��|w��-dp����#������ x���PhP�8ۢ��f�u5�eb'L�Us�o�[B�+�R��u��VM��i�y��+�
��#���Йȯ	�� ��E=s��(���a|��u�KG��L�����[]��+=I�`���4�N	�a�=?�o�U��u��ˁ�'X0�M�mX�.~\�d�1;�Z:*l�
U![�w��Y$�7rc:���+�&�Y�D�1��i�0��t�n�q�˸,]P��6⌥��K��� xA��@�S��aXT'��8���l���9v�Ĵ�{�:��U�w:���j�GS��)�CV���1�r_U���Im�y��Pf����������<~;�Q��.1k�r��v���B�e^B!���T{5���\i�Zb!�G�q����t����l3�W�=�Y�$"��˹f�`qu �?Ed+��0L���1L.�f��O:e��t��%����d�(Ƭ{��$ﶰ=���=6�
Ŕ恜�������^E�W<��J`�2�K��:�Ս�o�[b:s�=�ف�O^3��B=:��&:�VyQLN���6��8t��_蕣�<:�fQ���@�j�G;MU��*,���XlxVHYEB    fa00    2a40္�.i)����YQ��5��<��~s�����ä�zt�+_��.���Ea��y@U�_�=�- �5FɷNU�2��l҂��	�0v�V�d����8��i�9��(��.�rE��^5��i;���E����I�T�c���D�W[�KW��L���d_�m�/&��sjF�[�s��U�������P\�������2���zEm#�������g.��>>�J�(~�x�Yre���;5O��X{���_��oŀ�kvg?ї@����v���F�=lJ��:!���!?��j�-�4��9j�a`�@12�?�OXp�G�0�1��od�7l�п��4���hP7u���FĲ�o�:
��:;z�ID��n�S'�2�f�X���̊�� �]��k��C��Ha~F�R���5P7�P�����˾e�0顈{�}��m7���a�x��g�ė3m�nÚuG�I�:��
:�����Eg��f��?���Lr�MrS(��Hct��ƕ�0�����������^�J�լլF�N']v�p&%�����Yv�;�К�(�9u��Xv�O�s'�h�w�B��(`�Aߦ�����0j�2>H�u1Fz���ؗ��e�gQ�7��Q�V���j�;�M��Vf0�rDe�����6��.�]ݧ�c�9��yW�$ǘ��k�*z��lZ�k�6{-a�I���ݲ-�<����K�A��}�{�ŅQ�P��;cX��-:����~]�$�R�\X�g������Z�}F"z���+�耢��HVf�5�̳E֑F<��!�I��C�z���G��g�t�ѿE�G&��8Τ`g�ɶ�4�%!�w�S��	^:s�|�|�?m�%Co\��~D���]t�$O�	��n$e[~8�����Xg�A�����w�.�HX#�#5"�P�Œ�?��0z`2�YE 7F��>�u��1�͹�053�8^x70�R�l�ݣ��_l���/d$F�J��)�J�\�!�׈�����B�k�v�����b*�5�<��Q�������K��Jr�˪��@����6�&:J��-��8���5^TnNa)J���ؓ��%0�cr,#�G�HF���]V�m�¬u�? {��[�칗�w��egS��B�t�$�L>�k^��]��c������Rf0�J�K�Wq�嶆�G��pD��%�A�gy�>�hL��g2<}CTDwD
���S���NM��P9���BcK�+�EЃ쇽���i�6(���5/��m*��h	�=U۟��,�s�.���(��l� r���kq���׳Hfb��oqMYX�0�����ד�t���L�[F\ar�D��@�WK����r|�������/W�ϔv��,m�����.��_.j��Ӡx��g6[�[�m�xO��*ʉ�-����L�����e�ϫcH����#ʑ��lg��L�~7lX���(*��W�hM��Ul$�\�́ߪԕV�;eh�qP8S�;'j�Z�	��5^	m(�)n����� M�k�,�D��"�8y86R㼟Z�e�,�G���:\��@��P����&��ib��b�9�<'e����q8d�ͤ��� ��?Q�*?O��͵3o�s�|�Iڕ�M[��ֺ��/6�S�Ț(�q\�^3���i��.�|ke�%��}����z~߫��q���Q����0ܽ���v��[U5`�e~�6;�k{��u���A"�W�@7/~H�+�$ D���������D,��B�nߔ�����;���Z�\J��G��&�bJ��g�Ө��r�N�OeͭdQ��*�
��3���`�8���T�W'�Ĥ����y"��!c#���hJ��N����Yu�5�+n>f��N���>����@���^�'|F͏��`k�����T1PW�Cn��H�����ڪO;����B�9�wI���Z�K�!d*Y�lf�mD���`��rI�����|W�B]G��=
�5�E0q{�ê3E*�v4�l��WغA�����&>b����x�n�����;�Nc��ٻk��� DԀɤ����`3l���-h?�L�4KM��
7o��<��b~MО� ~�ͻ��+1�-��HM/ Wj�E�:GP��
�ͯ�O��nN�?X�5�J�.y�`m����Q�����<N��f]n ��צ���]a$�e���Q�c$�q�_)û2��&c��ǯ���2�t�U�Ջg��ٖ����[P����J�s����ѭt��U5��.�)�|/gN�3y>)|y�!wi�E��W<���W�F��祁"�C<��ِD��/!pŅ;�pG�'�Ƴ"�p�Ԝ�=#b���	�*�c����JT�<����܉z���$�囷
�����:UŁ\��,ų����;`��;KZ;���]ö�9P:+K���Ԅ�)A�UL!%�mk��`i�û��yo�Ӣ<����;@_�ow���p��u����뺍V����I��#��Ün��7�ӆN�Z;N3M�8�̮*'����%ׂMB0�#<�L��.�(�U"�M�k�3��+�!�<��-��oJ�=��i��4�g�4B&�v<��s�>Q3����0F�XO6D�'�:��N⿌�]��6��N����=h;d,:�1i����� {�pO��*�謺`F�u��'�Q#;w����-ߝ]�#�?�ˊC@%	�9v��U*��������$��:�����v�ked����p.��k`
�̒r�-�������m�����]�eq�"��+�b"4 ;�}����؇�4Ha聬���{�PH`/�=)���Ӊ)�w`-\��O��<�3e����EK�2������	�T��+1l��VJ��{�l��o;j�It�E[�	{5Su~?�+_7U��u�^	�;uB-Ɠ��#""��
�;C-���yU�X�DY�檯�Q��4��`��wڂ�� ��Q`�_����t���;oO�?V������gV�Ɗ�q#_+pQ��d����	���u��[���HY��G�C; uBV�~�-0�/��#�wH��ә��xv�&�&B��L�!��	��d�y�OmR�O�������	�c�
��5��m
ooc�����e�t����T��W����D�?C�vR`+j��:�#����H�R%����;p�{�J`.���5?��l x��2���M��07��9=��#�χ��3w�2R�iiu�!��s@�(��gܭ�����e8�B��@�|�H��$��Jȋx�ƻ4��V��Q���@�T��I|Ӳ�c���X��*y�_���7�{8C�|�������29�
��|v��'����vBH��%͐"�c�DF_V��X$�D�����e�\ۃ�.�|F�y듅�}�'*h��{V)��iW�.����w�aW&*�W�Jھ�h�=&Iw�5�
tE3� ���Q|k����o�2&xD��]/�P\�N�Gf��n��qj��6H�VY{{��;Ŀ�밶���D���@[a�����N�N�?�;�HK�L �)�'��a�VE{H�x�
�l�Կ���z�I2������?L��_������DF��x'�Y�Өv��tr�©�b���W��Rt;����@H�j5@֥�B��*���9����>��
LF�"���N������;Õoh�A��x�{�Z�a��s�5����'�J���߽;!�I{�qUI�KJ�F�3���08o㿦���4 8�����_0�e���Ȝ���#�TU܋{%'�u�B7�V��Y���`µ���+�S�JA"���}V�Z:۰�i ����R~/@�+�?;�7c����"��}eW+��C��HO]���L��f(-��Oq��'��'sm�Z���E�x�gG�������\]�݁'�'�`���~��t<x�3#�hM�ɍj����8��*N[��f�wm��{m�G:z�>Qخ#I��x��{��4����`� 3�ɵV%��C��Q9k�U�k�3±���H���p��6��ڭz.��~qi�L
� �:O���~)Tg{��4�qde�C�<�(���^���&_�R-�I��]�}��i��	&�uK�G8�С�iU��4�"��Hn��`�+V�T�(�%���&>?�= 0��� �%�Ċ�=�KL�Uq��[6�%�O3?wa�)h%���{(qH��V��М������uAhu
�L�h#��H�g�L�^�mE�%?���S�yȽd��
R�pL��1�E��l���揬�X�H�y�cPNԝ��b$��nb:�6�BC��~���}�Z�13ˈ�,�_��D-��,w�4�)�1^�t�\S6��8r�����2�s�WcP��rŖg��4p]����j�D���j�h��O e�w��Q�8ҝN�n�Q�>m��)<J'�hVצ��㻀����X�f�*��П��[}�4�Ք��#�ey���H�n7�s� ?�L����+x-<�hؼ#]�*���+�\�NL;���6�b%��r~��^�AJf6B¡�����$��/��A�`��9���Ԏ���#��KR���5�L��|�X�e��4-��۬n���)�}o���]�G(l��m��U7,SsY��*�{5t��p5H�qʉ����^�Cf���ZN �1���R��;��7��h����
�#�K��5����tD���^-,��f���(�h��o
��HSIeTӥ���F_���t�1��jJ<���~2� 2���=��P��� I��.fZ�^\������f�jm�,�2r�d�d/G��ECo��V�ì�\t�kS�Vޡ�	�hM�BR�ߛk�=t�=���!~��e;��h�dyYC�IQ�*e������k�S4V�U_~9t��{v��0��f2~�0��/x�����Bۇ�,�LvSW������}aa|h�"��(�uK���Q(	(L�V���֢^8�[�j��lLm"C���G���v�G�1xYOё��|�(��𕯡z�N�5�<W
X%�ʾ�"�R�+b�0+����v�
NQTSy�NȐ�D0����s��"
�eF5y��`7~����� ��:&gS�>f6I�!)��81?.j�����Z�	��>�x��h%�}j�?����Jh�K^�=�5 %,C��7i�Ѧ�Av��8�A1�˂�q�E"�,��QͿ#}|�ۋ�7��F�7Gz��-{~���l�9ˆX�|\J<�5UT6}CN�'�g�Cu��T�z��R�*�T�!��;�tt���@�<�A��-z�<��INe�a���k¬��\t���R�A*fB>kʷ�A��;0�P��/�K��������s��y��pr��+�rs%~�E��nV�Ό��߱W�!HW�3���-��Ѯ��q��Qo�gY2剄�dd��_}�u��@��ާ�X;q�=�\��ӄ	���,�M�� ��k�����k�C��xQ.�D�n�����<R��7ݼ�b��dlZ�g�.��
G���<	J��@��md��9��4P|�ƶƁ�H��>6"e � �(
���k^Ykp�ו^r�[m}؅.�7��~npqX�5����n}Z���~Btɾv��\���L4���S��43�+�¿��Ez�17<*�.]8��m�O�եN{�m�: p�zT�EH`��bm<x��F�?��>���$��x�����f۞3���y��Ϗ�н��V��Z:�� �1� �0ߛ>���K��f����ҷ�1���^1�/���W/zx��~�~�ſ�h��o�K]�ڨ�{�i�|�<�,�à��Q�0�+�B��noTL�������?�
B���F��7��H�Z/��������gi��!V�� �`Qp�gձ#t<vy̜�,���F\Ȃc%xMS����Ȏ!�
&Z�;��AU�ެa#| y��#���2MxiQ�s;��l��c�Jg��?�w��"Lm�mhK?�w��F���{.�η�����бv�S}T{#�m���k�l7�'G�3�e{��gP���%�[$�=2g�K�A��a���p��-�@uR��x`������/ghW����]��G�)�]*,��T�����| LHkܤ���G%0�rds�iG����Sk h�ɑ�?ܰ'Mw5
W 6!��w�֗�kw��L��b,u�IXe�+�QT�� ���C|�e�T������3�w�og������OU�@���]�_�;}�� )����[����.mq��J	xQwJ]8�X)e�b0�ˑ�L.�j�	��&D����;k,J�.z��K1�����nm`��Q`5���^ �G�w�[���U��'�S#�������	�pr���RJ�4l��'{8�~	�>�M[��z;������#�ko��xѴ����Ϡ�Rؼ~0Ư10�[4ie��Z�V���f%��垿���n*xUd�Y=�^�����HH��_GZB�+*�܅5�"��@�M��-J�UTU� ��t��`�ʹVZX�MGyT�er̫���3%�����4���|��"t�GŠh�]RЬ%F�e9��,1����I���=��C�,�h�f��J%[&'h#���0��<ƽ[H�����+8&u��Zz��(%�����q�x��Z��?Q�|;�z�P3ĪLj�]��DA����mW�i���m��*8��"�-͜B>b~ο�����Kd}NE*іjϱ��vP��O�^������{ǎ�0sib�m�ȈU@�րS��^؋`������b��^��T��Hj�fE����[��0��!���ǩ����u�%TP�k	O%Ɨ�zq@4&�^ly�@	��7��B�,#�Ce`�����O�/�?������8=�s,V*�6ZcB�x�6X� ���U����͗9w��Zt�v�͐��,���zT�5��@M<��{Й��/����C̡(�ȇN�;�Ю�F���t��z!���%M0�#~;O���{�@ݟK���`"��΁�r����#�,�R嚴�XR�<����D|�aț��M������m��$��s_!!Atj����?���G�C��l���)G:�1�E�+��g���\���({���q�Y�؜.a(c>_��S���R-t�������?iZ��Ůz�I�f7��MgҝF��$	��W1F�M�3�s�`�x��f������'��C+��}O�Q�e�=��a��vp��\�Q��;o����,����ۀ�!��u��oo��IÍ׷�`�_������R���Z��L�NK����]z\c�C�B�[\j��$v1�Xs�S����v�?�^���̔��O��\�]/���v�4(��n)�}�J�sC�ٗ��⸌_튥�m]bĐ�D��Fn;]�g�i�7��;��!�h��Z�IX��\
U��Lv��cJ�7��w�I �!DbVs�`���h�&�=����.8�&��X��j*j0&��b��p[qΈ���_�g�����a�.���<������ X+T7�(r+*�*�ec람H[��Q��b�Fx>�q���7=j�y��ݳ@�$�~Н
��9���	��FY�(䗊%�]�� 5���*4�}~�f��_R�-vz׃ނ�́�.��d[MUY�%�~�#/��\0�
��-?���AD҅���Vr������Q*G�d(����wק����U7�ʤ��2#yD�[�}���S�,�hA�e$s�ab}��n�̗�2w� ���m���F�1��Q�9zj�6~��UM���y���\�b��v��s+���@�ݤ���� X і���Ș���b��~�a,�[��*�q��f��)�:�aɅK��Z���E����^�[#dW��g#k<�{� �)	���}�ɞm�o_j@�;��;	~ύҬ�$;�fsX�OO�a"FG�7�Jݼ/�c�ͧ�@%�|�u6�L��>8�ʊ��f�S�׸��ix�5�٨t���8ve..��[��7�4�Hnj&J�/a�Ϙ�B�xL��:p��T�K <ٸ�X݌�L/�P�� �M���ֱܛ��~09����������za -�Ѧ�u�9%�ɟ�4�O��Z���ER�����֤�MLe:^@�Tc��<j��Hkj��<kn7\�*CC������Mu��:-��
���)��n�5�K_0��2�n��w���И�5 �S��L-(�o��`Zs��2��Ҷ g�{��"_�Ϻ�dhY�ǯ�+�.���G� �Ǹ��K�#�e
ƍ
��)��$���M� ���c������3�����Δ���|çG�q�7Tϔ�x�^$eS��E�H1l�K{!�ޭ�qΒd �6�O�Z�N$�%�.5*sL�0�1�5dz����:�lƯ��A؏\�Ǆ�� ��}ɍ�~�-2�/�p���q�UhỎ4��sL|'/�J�d�������G�𼄼�V�d~��:j�O�UjR��i5hMVْ�=E�W�<\p��Tv���Ed%�G��5~��_�m�ޱ�0���_�����iA���.���6/ �����3�ɜ���;� +��(���>>qb�+���Ⱦ4I�&=�7V���UUv���)E�I�+��|eH�}�����U�����ً����Dq��1�����B�=��(���4��T$A�E�����T@��DB&����3Ӻ\ق�	�B�4�U�I��7�!�cM�Q��a�j!�n��S�i�R*�Y��:t6P4w��$̏�־�Ȋ�Sp�BVP*=��t���.�V�A�_��G��A����0n���?A嬁IVD�d'� ��&�,�&�o�#X��(:�@��h�р��	ɬ8Ű��(Y�l��i�Ii��sq˂&Z"��ҁTt�{u����~>|�?��T�4�5W���D���\-~�z��S��g;�ez��]�6���.�@��̑)��5�Mg:��2�U�ᯕ��'�a�*���;+�\b'��z��x�vںtFu�O�O�i��� ��&)ӆ��<����/��٭�?�8S��>�#�N	ܤ���&2$�c{HNެ$�.�`h'Ҁ��z,]�G����[�ꢑ���E��-I���n��&�O����Z*�M�Ȑ,��@?V!J�=��Frp��X�bD��U����[]�J��v�l�|2R[|���5��:�H#f'��7�$k�$pp���;����IYU�9믙�.�l�u����'�av�Jr=԰��k�Bˉ�h�TY34_�*œ�x�أYMi/x �}z��z�~�.@�@��������e}��������E���AmZ�����E
'	�T���1���Vܨ��@�[��� 8 :Ăb[��!:��w2a
�N��ݜc�'��n�&�������֏L����ϐ/z�q��2���o'+=�-i�9yʐ��P�TnL�/�DZoi����R5i�vT�K*��}@����#��4�3�,���G�u6)s~k\ŞWа������2۱��Ɍ�I���c+t�-�-I� �E�� ���t>��Z�uFZ؄o�m�!$�(7�;*���d��^s� W��*��H��d����?�H
T�|����1wנ���q8�Pu�+�C#;�c{櫝έ��R�{�l��V��y�r>A�,��'X)��'�e&����*	#����n�����h�K#`����X	����|�y%�yq�Zَ���V~�Dө�r0��cR9p�����r7��Q�ڐu�>E�e�ԌP~nFX�a�o/QY���onxNi�{;�d��ʂ��/��b��T��������";*ŝ?��|i�S:sf.uEa��۸$�����A���
�9(̇�w��J�ʰ ��e3�l-M� �lpUaY6@�{�E&�_s	�Q�C���L-u�
�X��!����s��4��Ï�!a��  ��������-����ⰄH�ks>���@�wOH�x�^@b{Q~6�Z�����勃`4~���r�ѧ�iPS�j�+ݒͅ�=`c����� Jm�A_BڀL�Z �EQ�A>X�2�K�Cf:��]�^	�u��)��*D�r�G���t�-#���5p��N��� f<1?���d���YЂ;bSa��3��a����[�h*��AC�����G�A4P���,0��i�l������~=ې\�+i��A����o�$��kb��a\�ӷ|?-�PZz���˪��Q��ʿ�,¿�M�O�+ҧ�h}%-�~�ds��P��IX� �6�ݍX��j�������YM1���n1��<5}L}� �tt�V ����n�C� m�Y���m��e��X�A�Ѥ뾨��qk:�1�)�MM�mɓ�p8fio�G�@y]a�ħ�h׺��ښPv��ٝ��K��
�e�~�Gr	Z���8K|08B�E�Y��"�*�D����m<%x>ODQ��
��O�(��z����!�	w��h�M�lʟ�#HB襣��Z�D���)����oܒQ� �����B�&�^v����Jr��V��2�>&�KmO�I SO0���98by�QG|6��3���v�C�.m��CE��3B��c#�n��QVm�'�R�(�NR�Gz�zMc�<	�u���>Xߨ������XlxVHYEB    fa00     8e06�#Q1S9"��"7�
��7�k��#Ĥ�	��a �5��h4Cs�u���+��t�j0���i���FJZ��'��-��.<�{غ�C�Y�{G��c`�0��o�W�<\�5?^�^;q��Y�(Z�Uq���=�����$��w��R���k�5�'� ���i�.�qO�0m��Ȉ't��$� Ԗg�~lC���T�&gA4���g=��*�;
0�g�S���8�m���Z���H(>:������TU̣z�Q!(픐{��6"v]c�mg�s����upcO��qg�R}^ҙ:)?a {�T�d���q>J�_j�}���_��l�ȝ�[�)D.I+N��?�ĩ�ܥ)�>�����/'L=G��$ �
�G�D5�����s�%��R����?B2��@�<��d+�B�G�����D]�;h2���in|+CmW�Tu����+��(�	7v�UzKw�ۗ���v2�Q�9nt�Mm�F�B@��<.*�e$n�v�ג)=宅�{i�BՄI�|$�v�^c�+�F�E�l�����S~)��F'��VI�.65�l#TV�E���2�܀Ek���s�r{�[<�9m�5+t�ܜ�&�R.ObL
�E?c�ϔ��]�l<L����; ���6x�̐��Fд�0NB(4�F�i�n�5c�ehVhL&����Ո�V�,� ��Y��ՋI�9�`�J
-��Y��/�O_dE�6	�p���jK䲰�5�^G�fl82�f�o�����G޸��v�8��Z��L��ٮ��v����A�)��L�,�=�������}��{�,�T��;�������%�{C��HhE�~�kE�8��܌�uÛ"\�9�J�a�+ew\���~��5?F����e?�SQ�.*��c�q9N�Q����>���?gģ�)��t|�?�w������e���!�@��zɀm��6��dI_�)�VSNE>:��p�Q^C��tX���������ZV���	�#�P��Ϋ}���N�R����ϕ���� +s��<z���k+%�0ۺV�U�AQ��"� L^��SYf�U���:��e�gi�p���z�^� ��Hb�@�����?]ᛐ�U�}��x����8��Z?��v��W�^�U�ht��1���R�Q̛-^UA�#������ێS����<�0�\�˴*m���c�+�ᒖ��Pd�P�e�{	��Ͱ���V�29X�PU�j����F1�ۦ��UnF�m碕ro��o?>0�����?w���WGIb��k�Pc�,����v�:ۇ��2V��]�
ԄiN�:Q e���Rn.�Th�_2΋��7G5w�F�5��d��oݕ%��r=��\"��ຬ^>%Fව J���m�����;j�=ӯ ���J��q��g����w�N��d���g
kzX5�yd��->��-�D��A�c&&'�TU�:	tDG��o� �d��&�O�6O����\�9`(8F:g��1Ku��@���:x�� �i.J 	a;��P ���n�;O�m�3�"�G�#�	u�4���5�{�VOV��wG��{'�MJ][ocL�:��dbd�f�sCR	�Տy{/����ı���i E^R�0�jJ����q���Г����:P8b2�^�\zO���خ�[��T�`��'�� �P��;����և -����O4k�,mՓ�v=�5VS�p���	�T���'̾��Ύ,0�<Z���ےՉ*���n$R��/���W_/�R�ǻv�:F�p�\F.�(�l/�X���*����M*Щ(5w�.9�{l�����sC�]�;���'��[���N�fd?�3���0���ڥ�'�s2�A���Tz�ƾ�vlow+�F�5+��V<B�瞈Y< k��l����w��I)BiY��K��I����eJx��ԑd;[m����
��viT��o�Tχ4��{_C���O_�k���ﾠ��X��0{|����>r}^�iVPw��ll�65Ԃ���Q�}܏c`��9Vhvm�[��P5:曬��sl d��ǽ�'�L;��4Z�ӭx�u��n���q8�����W���!ѧ��ÉDS�L�����6T�5�]g�,�X��[_�	�>'e�A��-����]Q�f��#Q�������O45v�qQ��լdtŮ\0�b�`R�*�ә/��bQ8n��kF�T4ğ^?fz�� Z3U�歍����T�XlxVHYEB    fa00    1110��Y�-{�ݣc�u%ʃ�C�>�B���uc�����+�=�1IO/�ky�$��N���+#zǨ�)B�Į������r��s2��A|B�p��r@c��� �1��};Yy�tmλ\�Y��x@�?���R��롉q����]�n�����*����d##��7��)�VH.�>M�r�w�'��k�F��q�Ѧ���= p���į'��8����!=Rk�dHԃ�{��Wko���M��Z��)�I����֝A����,`K;���=Y���������S�1s���l�8��uG��!h���!�O��:;c�84�A��ṹ�6�j�����4ѫo[!KE�!���PㄋҶ�J���3�2�j�J��0�?�&As��Ւ�u����ޔk,���E|�jnvJU�OVuG�R�D/�p̻}�F���i��t���z�T:$q�mF�_B:C���)��xPa�kL�ϸ��{�K�/x/��xE��]a�Ĩ�*�w̠�j����7����W����7�6�#2���5�nƓ_���ܷ0	C8x@� �V�i�A5^_�����~|�
����C[�}�A�Z�%N�u�\����X<�.&/���d�*�r ��f��JTY� u�i�����V���"�3x��G���f�$ױG��A�zN�%L&�>��C]�A�mzە��!����`�\��܏J�"I�ǩ�_��p�PH��D�Ai�K�)[�	�0���$!�s՚�Z�.�������m�-7��1��Λ6�x���?6�H���#��m����R����r�h�-����-����X�k�X��6S��%\+ґP�S	�%�8#䞻�/,� ���aG�o�M�Ĩ����$�n)3&��,�K��Fw���������Km�H5�����Z	ށh���C.���l��AZ����-��T9�.����	H�,$��������54�j�@H $���P�a��5O�_��x�k[����:��x^BẎ�������rXmN���:zi����AC_�t�'�u���H	�e(q+���9"�!u�E����|�)��u'�)�z%H��{��ú�������Wt��9�Qr$�5�'�Iö6}�*�51�O�.Ȥh%ّ��,��2����)<P��uN��?֌����J��<]�OU0�$-��]?��&-QA� Xs3��/Rf�:��! :�6���_S����9�[��%�3~��s�3��֏�k�?�r��(�����~<S&���X�2wB�fD)��X\���u�>���
v��JՁ��,�����m��УD�SnDa���L�CV���D8۱�0�WMh���n�}�	���ٺ��KA�X����5|Z2�Mi]�K����2숶�h�\R�TS�����w��Q��OKt�a<�؜+���BO�۾����"Y�~����o������ІF�
�Tv&�x�#�Ѹ������o[�N1G��6��ke;�2��^��*(�}��>�S0`�����W�����b��V�`�3*�=z�[^y=9��dm`f���r�"�i��GG�;i��F&�t�l�6�����3��<o�����޳1�ډ���9� �_M�2<���]������+��L���h�~�G�*x#��m�t(�<�yU���ےz������}?�>�P�Z�F�'�9Q��8�� (�����G��zG����f�Me'�}�6�V�l��p����AZ3�n�D�OqT[5�e凌a9���Q�/Y�̋��3�c	�qr��˅<�\. �B�_W�i�bE�\�NG�o�㲸�r�GRU/~���>��.hQ��Hp���2(�R��f�i����y��*;]��0��	��H�F�9�W�O��bk4.2��^]O��>���E�o<��:pǐK�v��M^��,�Fd����V����5��Ct��Q�`�<_�B<Ø>"L=���>F��_cHĴ�j���\C���Zy�����|�a��WX�'�	�E�V�u�<�%�M��;��>܁�\�1��j��%I�(��sG���/C�ffV���M��d�$WQ�1W(��C���K�QZ�{Л�E=�~3�r� g��<��>mi����D�=��*A,1 �ey�_J�zq��9�������Ŀh�E��/lҌ��XT�B���R��d�*��G�X�9�T�j��QD�-�2���d��ktI�<�s�'�t�~�["1���#JbH-�]�
t�n��X��>�?]���A��4R5�W�jo���ý��-Kԣ�&�S)���x@�Ve�ַ�b_.Q��1*� GĪv��kF}0-�:%��@Tr�7�L�d�t���Ν�������+�3�����Y�C�|k�q�nQ�_-�-<d�P�w�F���-�E%\�J�[윒�4O'��g	ۣ�+(@���v~���:���[�M:�;5�9�i<�ꙡ���j5��	��$�ı�������T��3JOm�}򺯗̕ ����� <HS�Y�9r���T���	�LZO[���$���J�;�}��9f��:�Ն	:� �+�'��\�
�ck��f�x�s-����i�����Z*N��늻�>���s�/���x����҂GA(k�ƐV@&�H��_ZS�.�j�3���,.
:���a"*����=���^a�e�2}�hwË^��N���"���AS�[p�>K:���*m}���/h�rxu���$�L�#�H@�݆{��?m�MHS%��ܩ���Q��Obi�)X�{B�p�]��eT(1�>n?Zb�f�Ao
8>o���0E:���� ��:�=˜�hጯ��G~o��w2��[��x]Σ��L�l��p�7�G��~$� b�#�M�d��!Nth�'���L#8�Ղ��,�*N�0�v���7W�O�%���f��i�\-��V��O��3|WV�;t��r���vM��P���������?kKYE�ŏݮ3��'S�ٺ����5�lT-$}�P�Y��{��0!��Ci!��1�ix�^����d���n�a;���_��y��*�����X����x�g����3~>�+�Gkcd��QM3�>.��p18�XD˺HMbk^v��seE@U� �H-��j�uu&K�|�J�v0�� ������lPC.�
�،w��q��b^t��#�W����R[��K�?0>q�(� "�!�J+͏S����'^6~�	_fc"�P�\��	��H��_9�"��C���ׇ(dm(�w���۹2&��;	$b��E�޴YY��`���mV����;z�{�k�n=+��g�ܭ}�-��A�)������vjI�7Z-Nz�6_`ՁI��`�;"LL]d�/��X�ʿ_�l'�g
�>����sVx^1��SZ��n*q]���p���S�eR�M��<��e4%���1��A{��V�y���p�n����~Bt���	�Aw����p�'<t_��0�|�{�C�&}�)<~`���GPӦ��=�AE��r�) /7�^0{Go�Յd�H-GEG���M.	^�9�o4�vw�YDǒ+�����ռ!�$���l�~S���˭
�F�*��s�ȓ���0Pg��*.�0��K2�`;��aǘ����x_��
H�����Xƌ&JB��^ޫp��k��=�qH�v�C�,�W����U׊����K�e��ɻ�>�m*�syc%`�v�$~gQ�AWۧA/�Yw��8_�-`$�%�$�b2��(&��Wb3���C �eg��[���pBt&TR������T�X�,�O���G�����M�Jm		�-*�nj��{F��R�z�y=�>����~U�*�|�`-��2�YsM�v�U`�j�s��J/�rZ�O&�B;oxRR��ef�l�K���</�y������r���P��Λ2=�R!��%/�~)�i8
l��5D���C?zO*"�(zS�?ȿ$�N^�]��!�?;�Ψ�l�(l�G05�����T&�t�逞�J����I}���/l�"	'?� ������Ύ^q?Ra�c~H��v�f�X+��j?���1���>q��2�(� ��H�7`����8T�������/�l��/یɴw��]�ǹ���S&��8�Q�	L����$�
�}��؁V��.��D���(a������&B5�lW�'�=(�������������	r��	�fa�0��T��`�~&K�mEVE�h��!7�"�5;r�+Km��@XlxVHYEB    fa00     ca06�����C��r��ym�C �b��P9)b�l��h�e8h�l/�!�A��yB���,#��Ft��s(�.5O��:TU g"Z4K�᧥n�m��.2>u�k��Y>d�ɛ8�k�P��Ď���وW�,����d�����*��W��VS	�@j&�y���˱A(,p�Y�T��8�1�z��KiK����L2����m����d147?> ��Xe}�B���@n̩R�B@�:G�^�k��o9��)SbV-�����<ұ�I��$�7�������M��О�sa��*wZ=$#J��d^DA�I6��k�$�Eg��z~1�MNV�
��/d9aʅ�_x�q��	�GVo1����_���V>���}���bL��up��v6:�t|[T��E(�ć_)�jn7`��@�%�]���8��m�ZcQ�b�4�O�L�J0J�(8=�\bU����R�{[��b���m��4�� F{�F��g��	[�~�׷�?�X1����9itnB� |x��0���m�ͭ�~�M����T+��QK�nP�-薨[����1��P*��ay��9`Guh�/�nS#_s�g�/��RɽJcS%�_�W�=1U���q�8��ՀҮ��k�Pu��Sį��7=�3(��Wƨ��I$���ۿ�c�s7��7X�9	}��Ф��B��FxK�G|�1�vs�K���z��C��RY0�L����wM�US,��a��w��[�"d[JxH��_��]L^Ԝ����{];j\�VO.���8��[��'&SgX��?�4�.RC���ǈ����p�p��;�J?yq�Z\ב�Bz�M�RT�J��wػn���t�2V�UQ��ܢ��.���YŖ�~:1쟸���H��:�� kq��^��2����ꈘ�(rȵ*UH��/�8�k�A�clC�����h~�Ъ�SS�F����ȑ�c?ߧƌ�Zol�?�)�5[���n�pu2����}f��h���4:j��q�p��B)�&�c�+�����'��;<�ˇ��FN�Σ�>W=qS�t���-��'�~&Uu�`�kx��ʢP,C���@ł0�\A��/s%��aS��g�D�%RV�נ�m��ў+0��/F�q�
l����F��9��,]�Ϊ���2�B���9AF������>	��$����2�L.y�C�M�=(R���	Xo�:��*�4�,�)q�2_���fIX��'�°�[onu4Ę��)��4���ѷ������nt|�H��� Z��ۋ�eI����W�kᕕ�5�@�B+�}y��>�Ho�ENX�^���㤻6������N�d����� ϑc$�5�!`��vy��1�W&�*�����#]a�{c*P�N��r���'����^gYBZ*�)���b@E���9��~��_�P�C�V��Z3�Q�m���TѺ�V��`���|�G9^��V��8ڱ�o�����8@w���p��b�z3�p�$�&��>�)�ܖ�N��sŮ
w�m�N���x*�e���o�<��@qд��C�͗v�Hީ3�a�_>5�g�@�耚9����6wؕ����t��6�׀DHs��~��TZ�b'^������Tf���� (�`��}��č�O�i��#��x��Ij$ ��wKgl��·���P�� �F���p�L�%�ߪ���Gj>EW��vN��I-	����)��D�7��m-$���>�,�������� ��c��l\ ��5�&ּ��;���-��\������X��N>8vm�}^0o(;�C�*8ޜ���lЕ��t�)�&�����}�B��G-sI\�MZrG������Ui"(�#hB��G��EA��*��h�����E/@���l�SV���E7�;�mcJj�g�M+��^l=�ɡF0���_�ؿ&:�)R>Rr���)�븎!�-'*��j����|��~Q�p�ȸ�C�w���rوHR�>c���f��[8���&9X���Pvr�PYԭ�i��@��)^�r��E�A��v�'*�/]J�7�pWy}"f�����+�Qt��Ͼ-C���w1Y�h�����<��<-EoQN�e���ӝ4��ObH��V�&�Hs���dƲ�e7�ߊH�]�]��}}�1�b�/\[��#�E�jčOI`����	�Q�_+�`���l	�h��qnd�ر��s���i�8W�׬�7�vEy��I!�[P���63�sQ���b��i횅\r�!m���B6Ce�Y�s���&V��&,
3��"�λ��iW ��f���yۅ�4M��$~�"�=�=�-�M]ow�ɬ��xj���K��z��.<̉� � qUj&�"�:e��s�Bv�s�Y��e���w�Q�CG�5��L�@De���ײ�X廷놚:�2�Ҧ_!���'�S\�1S�Ky6�Z6���2,��jp�G
V�ܼVk;��Ih�$Z�q"h�Y�{;5j��R�xl�$�oj�L7ǌ���,�=/��rCZ1~4���L�3��z�Ց�h�Ԁ�wO�>#b�M�
�iH֝h��]/�y�Ѡ}E��P=mQ��c�"-��Z~����8
��~`�	Q�����j�+���}z�8�[�K����,���gE��j�\Ր�j�ܚ�p�f�D����	`���P�7@��R�`�K�I�t�Yg����~��Wqo���-耬�d�L5��wX'���FJ#�xK_���|��z
v�s��q372�H�=�ua8��Vb���k�B��c�:�p|��=\ru�h��.� �0N�Jإ��Y����ߡ-^��MS>��P�OB�Zlߢ5u�0��Z���MUHyIH�qT�pK1�ǢSnu�+
8^�N�X���ڛ=Œt'��B�*�,_hx��JV�'�n�T�՛��9(�v���:v��N�p���,u.� �xnm;D��}hC�{�P�%�&���Ki�\YVVl�%�G/�F��ʇl�r$����D����q ��O������Ϩ�cB.�K]�0�����Oi8Le$�)�O]%��F\]�G��I'_:�t��!A}}C%�"��;082RQe�eŴ��^oHr]t[�u~!�¾�M��4)!}�h�wc��t�� S�8��ۓa6�0�����o 8�F�I�_f�xJ*�7k�{��QjGͮ�9#���4XlxVHYEB    fa00     3f0֪��v� �.-������զ��������\=&�c����M�x���z p�-��)��l�Y��Պ���u����:�m3�ZV�����UW+W�|o�{�_�Zt��'���X�e�����]p� O80�����%��$|*��֚�܊S�ȥwY'�*�Xa��a�ҹ�3�o�0�Y���=-���0K�5�č���k"�c�<���"�Ѷ�0��,H&���m�~|�r��ףE>��ӌcQj{�ӂH�f
C�9� F���8��`����A�㺇d7s�'�3����4�DO`�����M1E_�٤�Ұ[-�q���c�8����@e�B��=��+R�D$B�'��i��dE�g��E�<���F�1?���O��t�l��z|1`�I�$:[ON�?�����j_B�^��5#�4q_>(af�b���FI řh>扬�I �R��s�b�I��a�ڒ��h�C�	�����8RI�ZK-U��_��͘�Js/�ZĪ�H]�2�Uo�FeF��9`�qW�]��!�<&Z��M���s#8eL���q$W:?�θ$#�p��:��
A�[�b��l��Z�O�ib��ZFCW.@zױ���o^KWh�o�dN=	Ι�\jAV~t>���z���5���
Ș�ݒ�E͘7rRI�E��/��]�i�B2�^DB��l����v��)9��!ڋ֠v������eC�<@JދI��ë&���/[Xz��&�7׽C���+p�d3C"*w�����p�;�;�%�c�LL`�=�"w�L�yg�n,l\%O��R�����/o��
����1
o,mA�'57��V;আ��:P%����)����;̹�HGXL�#�Ը�&R�� tѯdVT�` {�~�FT�sp
F`����W8E��f\?-M��r'�dHf�Аr:��+՛�F�)5?d-Ϻ�ޯ���V3��2��y8�U����\>i3*�c���8\žV��j�����>XlxVHYEB    8096     b20���?����Q=5���t�V.�G�/=Qb��R_���h���,JPW��L�2[H�g��T�~��.L45�g�S�E5&;�/;H0���E�C'�ewJ�h��*�]/�v�bВ�3�Bx��Ś�:II�B4=�*¼�a4P˶�aZb���ؗ�7O�oK�0�;c�l"�|U�t�I�oѹ6t�5B1��Of>�hZ� gz�N�cx]�9G�C���C� e2���ݽ��;�I��O��#�B���Ҍ���-���9	������QQS.��9Pp%�y�Z���B���h
��AA��s�PPj�p�^�ϱ�xa��I2��%�P����D��QE�a��hnj��Xo�΁%��^�(o���E��o�Od{�d��{�kf��Gb�����,�(rF|����oņ���n��{�:�S��(�!/���K���T��}�]Z�V���(��·�|Z����{��Nv���Ty��k̘�Hp�d��g�-��|���b��C�Z�f�-�����"����E���i�X)��������bHJW�߯�ϔ4�ҚF+����&*�7��
/O�����M{Mt��3��׆i:*��CrB��7nq�	0pj���j�~�n�㿼��[*���@|^�ޞ��(xإ�k�kJ�o���Qb��a��z�i�rT������KL
a�L�
��nф�u��!�$��-�Q
�fI�1/�RK�@k�+���sS�X{��m���pi_�Q������M�η�5/�h�t`g ��� ��5X���l�<�c.�<��Syd�/}t�q��r�J��-,��NJA_<@��d�M*���
|�5u���Qڵ�� [7��Q��;PlP��x� ��`��c�^�	`��ń.4�N��h����6�ݣ�E��HB��>#����j�����.�
����q��=Q� JH��~�O��h@qp�\����vGF���j�l6�T���.�}������S3����@���R9��x8XB����ħȄ��H�_H�g2�Q2�V����Z�K_�.{���u88�P0�}�k�k�v� ��E����;���Iބ�<�޼xݭ}��MF_���Җ������y�
BD�0��Ȅ1�a������Rn	O��GR��?�����À�����)c��z�h�s@�hP&H��儂��*�y�ߡH�?�\��x���6�k�,������n�zq�]@"kّ��_
�$�Db(I�V�dƵsa���/�V��m�I�$�]����.�-f�h:�g�kP
v�����$b���|��5��fU[�5=�Rn�z?5���s�S�K�H�����?�g(����c�H�K��"�i��bQ�A?��ٺA����=ZHΨMǕ����S$1P����M�2T1���K(dur^�>��y�WZ�����2�f>��\�%�'.'=�?�+xޏ��`8ގ6w�J`��'�[sN*'�����*|���mZ��7���8\P�U��I���ft�ζ���/̛�*��,���
6$G(����bv��/��%t��s.t�%2����<`rPt��0D��5O�Vr]3��-gD6|��d�UX�?��|(Ws�A�����q��Rn�'�jL��	q�b���}ߢ����5|�#x�N�f�~|�]K����v�MY��zɊ4e�%�0�F����Sb�K�t�9iƢ��r���~���)���C{"��fO�3�'�o;#������%^$���Tb���s����Q4n����B�=C=��FȧE�p�sG�U"�p�.gEэ��F�_L������Zd|��\8OR�����7^�W�o�;a�]�q�D�����)�^23O�D#{��&$�^�M���o)d����{>QI�u��9~������~�]��ڭTe#?Mm6���{ö$ՔtB�������8(�P.�7����}�z�8�k��c�7N2��hUC��-�xќ�c|���8:J��Aa[�Ӣ̡)8��d�C@(Q	 ���&h$��g�o^܀������U�ETu��4f�1sA��l�l�&VI3tLM~�1�q��v�F?�8A���/����ܳ6��æ�#'�ޒ�a��dO~.�|���V�oq��eZ�U�D I֘~�-�C������)䩅O����MȒ�l
�b���t&;��/���gh��`m[`��^��Z���iԀb'��s|%�3?GZ׹��ܢUv�L��^3�胸�h�cV�~�J3�3�?p:VQ#+g���P�O�b�jxJ�er�a�4QÕ���E���Gt��x׹�+���n
�����Z�	�5����H��!Î]S�����<��������]n��(N��rwUP[�1	���	-X��>�Z�*��_ԍ���T�{\u�"h�W}~�C���3�d'��\���y�됗}`�|��,�7j�5$�Q���Q�)z�����X���-����6?D��c�
�&���ȏq�J��`�����g���ii~i��߅
�����W�f��H=�ʽL; ��� #��$P�%�l�LC�ea�nI���,�����c���}v�v/ι��iV���n��eE�8�	�-�9E5���08	>���k-OK�].y���D�C�,��i	>�	iF��,Om��d��
��ڹdń�[��E��x}��&�$���3����"}W���p�K���lOV��J&(����e�^�G�� H���6�m���>BȘ-�\�%U�����˛��q�Ŭs}L�?�tP�ӕ�ʺ�-u�G���C��v