XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�fau�'IX�Ñ��-��DZ�bރ���-���{Y��&/zOf3m%R�D�ǂ����B�fXZ�-�����%q7	�l�����7�#X�"}�W�sGFM�=E1=ɵ��a�h��`���\���M=��N4x���.�i���s���'��[������Oak����_�Ig�M
�*U),�c0pj��@��9k?���N8+{T���	��\x�C8�˔�SI4�;����q1ւ��y3�<�-1��|��j�E]:�P�j;�8*���������[���ά��f���H$��i��U�ُH`���D��]'���<5V�p1e9�C��cq<nrTF��g����a�*����u��!n��r�3GΘkŀł���������~����Ģ�r#L��u*��8�&��,�h!v�3� �� A��G(H��;�A�>�n#$�M\�����5���?+jb�M�/��`D��4�^C�fl%�+��t~�ϴw�wa��l[���]V�V����C��[��ء��&�����ۮ#�k_��Oh�o��kI9�Lm[�=���$µ���D<�lXR�Mȁra3k�hڈdx#Ҕ �N=�D�8Gl\Py���,1>yVD�O�)o�{,J��̈́�U����L�����Zp�Mu�<9d{.^�I�#K7aiK����?��~O�-�T|ca��*��pT�!pKey�c���|�҇�-�׾�'k��;��#cm�CQ���8JS��XlxVHYEB    fa00    2040͈O���t%�f\'����ts��צJ2ݑ`��7Dc��HG~p��f��f��Q�X�xm=
�?�T�zb�,x�)��i-���L�� �ִD��F�ǳ��LF�Ķ*b�=Ѽv5k�3�ǽ��kH#������(噓v�ْgeG��]�
hb8���������6'����Yړ(��`fc[%);&���e��>p���):���� !�W4�8��kz�z#�9�jN�;e���Z�`���!���8B�B��@dR�c/��A��߇"$Z�����m�@�][0P�A�iƚ�)œ��#N�*u��@h"`�Դ��ov�c��L
SK=8�+Wiru�4��R�p�9�HA`M2#Ť����J�=��PFw ^�\[�c��e|�a+�w ���S�(]�gY��y蕋���C��l�2G�@z����[S֖�����s�R�ӊ�j'f
X%�� �3�?�%pM�o=[>�(:�'�
f�D���:Y�"���p�oꈼ��(GB�'0b?y��D2n 5��聟Ƒ�:2BܒhBF���I
�ʣ
��{ݐ�C�r+)�H�]��A;Qa�Ҫ���)�����$	��v�x�V��ueYY! �S�V
�mv+\��IJ3��-�+�hIȿO��}��Β���2ʼH����#]���'�2D��_��>���C`���XG��ܼ?>����kRU�@x�#��u�TE����D��͕y,�SG,�zFÚ'Q����&w�a�hл!�z�=e��g,GML�q6�����[�!4���^���//AT�Ӌ�?M���U���^xgwK������vWɧV�gA���Y�E�"Z���Gv�UI��W��g��+G���W�v{Z����L��sm��eP�	I� �'�9�WZ�M�k��Z�:�gM�+�Q�����8�{�1��']C���*�q����m��S�Yp��P�F��J�	�xA�
�$nݲ��ȥ���� D�<G�Eɕ4j��3��A�� f�����H{�n��[�G%�C���5(���e&n �,�EA��?�~��E�f/z��gu��H�� ��i��J�e�>5Z�9즷.�F~� �k_�����_��5��]t��x��&�]O�jʹ�!��o
��F�hߦ�Μ��7P��\P�gi�ײ�����H�����w�����j�8�JX�\4�X7��&0�$���ҍmG�R�\�"��-A��� v
�p��mT���s=���~a�-�i��n:�W��>�=0 �(�D�,�>j_���k�Z85!�B5*J����_i���q������D ;�y=�*�:�����Y���+�������n�Q3I�X}�FQN����60P&MK�V�6��v�7����,�/HvH���肗d�l�,az;_�?�y;]O�}��z������Z������M�$��g�9�X�q�+'����toM��qK�e���CK�N��,AI�Iz�(k	|���fĪ�|m�c���禞k?S����R�n��4X-��-kn��ص�p�;���xl��:���ؐQ">�V=	7ýw�J�{��g ���b
)2 �\�X�M{d������/�#%���]NrS�zuN U�	�������I�Sm�N�{�*�
�1h�e���,
�"�Q��m'Qd2�lM��dU��ܟ���C_��a�n:$e�u&�?"��9Z��0�i���_�������\��[��
�#��I��:���+�'uɺ���z�e#�����O�	�P�pς5E�@�d��}I��SrS��rb��{s����ϒ��Lk��'�#�sP�]�}��>A`��3���I(aR�ő^�Gvdq�o8�v���P��;�{Bb:(�f_���)��V��^��,�E�&Z��xg��d�Y-�&cZ�!��"��DTA'�?�^d�����Н�@�^�`�ݔ~��5�b.}��?��m�97�z��=X��6\W���A��z&�S���cn?������Z�P�l0��vg��� G�oj ���2(7�^�} %�LE�{w������Ms�FTR��2Z���5_y���G	8)zN)F4���!����S�����y���,+�m���!vE�kzQ��~OpSH�Fl��KǱ��i�/�ȓH@��@?����?-=w1�q�Q�=v�E4�<��$��i+����Q����@�_���F��&��"�*���ULk��ۑ1*��O�
[��j	xrP��2	r��fn���f����>'C�n�A�+���.�`e�+/(%����t�Wrh���h ��V.'�i�9o�@�M�캎�,\߅�י(�4�1'%�C���1�K����E�8�s=��+<_��PA�a#6/��Rr�C7½��N
��>"�0��P86�p�Єԙ/�B��*/��#�X�`J��:����{xV^˒x-@��$*���%��et$�����S�j�s�P��s�nLq�
�*�~�H�-3-$7��d-���C[��UF.�!n�ʼe�G$��8�ʂ�ʱH�jRF�i;�d����Y3s�Γձ�'�0�lD�ϢxI3s�_b�����h6�_����`Dp��7�`��N�U�A�l�7Q�8(�M;|9mf�'EZO��P�
sD!�׭�D��a�R��p���q�*ܧ�^�����,��Ǩ���[�Ş{��l`�f腛ƍc*{n�X5���M'��p��(�6\�hR�"�?����{ۡ��l6r-;���OM���K���6������J��S^��GE����E�`�!�u�LC.#��/!1ї�")�WT����x��\��$��m�䉜�.�ǝ��y�N�̮c�^k�t`)ܫ�>�uA`7�
�p���Zň���ZK	1٨��0V�X�R�����~K��c0�}�Z�,�B�w��w�����z� à|��@�"�`X[:<.8���8��a (��'{��O�x�vu�ia����^�8N߻dgu�|ri�>��J�v-y����Ih�{�����U��o0{���b��ͮ�����F8 K��0�o��N�q�`�<�*1����B[�J�\]{骹�Au�fj(q���ɀO��Q#��ȡ�H��ۘ#�8��sҶq�z)�|�`�
BS���su��X�2d&z~��5%�9�z�ʓ!�?sn�:�M}����FSq-@ߛ `����@��5���|b����T7�>��푺�����;W��w��o� ʿ��`��̰o B�_tO�:;���@rE�����U�C��^+OZ��%M!�jfZ�~�]�9�P�h�dviF2�߉Qr#��p����DkLm��`�D�Ą#L<{�R��d�qװY���E��/��
�f-�����QO+�]�o��w�a~��ǟ��s�h�HD���{|�� ���"u�@�:�<m����to����II�6��¡Ђ��l��tٿ*���4�8WcBb��I�ږ�°
ڭdE���f,\�h����/��w������$���?����y�d��������O�F4f�Ǝkʼ�JP〈w�E����;,5�.ꢷ|c��W��9)�f�)����o0���m�+������=EٌJ/K��pz�Q���i��ۑ�ǖ�����QlT�\DQ?���O91���M�g��7�3�*�̣pNH��3h�ʦ�C>*��~HJm���G�Sw2:*r��y/5_�;�D�V�2]򣱁��gMK44��f��#���FCK�Sy���a��ơ��Ny�9[�TQg*x%,��7��N<B�Fp\0�31U�K?�rA]�bҒ^�B������-~�t�H�yu��g>��֐Q�x�h�"pj8G�y��A�����􏒑��$M݈��f�g�R_jv^�j�������\-����kM|��.�!��%/�H��[�����L������w�`��_�$ɝ�d�\C�=-T=�O��nyΈ���Y.f����:��$��YUj�f& Cc���~���hR�=�-(���x�����jnǢ��+�4?�vW�������M�s�/�?�#���@� ���;��.覙��>G<m�hW0)Zؕ�����9��;��*��h��iWn�J!�1%�2g��|�H��aU?"S{�2��W���Gߤj�=\53g,�4�EG��J����M9��Ί��ZQ�J������ջ�3���,
��X�yy}l���H����������_E�.�.O���E�
8��&���2��4���锄��E�*�۪�,z�Ѹbm�ֻ�x��0}Vng\+�@>3��2Y���F-[��U����	��+���X�|I�m]?P:��q�O���*jix����u)w\�d���s�I�;	@�o=��)9i':����/<z��^�4Cٛ\�*Γ��>h��z�b��a�{��X�O�9��$k�8Y��0ߪa��L�� <�QO��A�ߣ��	��%T~sAQj� ����A�f=�l��i��0�B�p]Ǎ�Q�"����!'�CJV�0����u�2!z��8=`h����J�/��VgI�~}h���IÀ��>����()~�����S�E�7ݶ)�E�BnF#�y�t��t�Vj��x&�2;�LƝ�uE��E�
)��Fr����32uDԄ��ѵ��r:*���'�?}��:`�R��PT|���	�w�����[s��p��#�´���R9P�$�I\�kXcgog�ڬT�k?�x���(]Ϳ_+l��w%g��Y����=��<���,cd�梳�:�z��c�� YO�s�@ra�k��l����hU�~c�n�~�Q~���;5�3rlӗ�N�@�����=�Զe��W��*���B���v�۫���n�=��uW����<_w�3xX��s?��� ���̌ɂ�����Bjw�3�Bxn���$��*�冃z�h�®F<�	+gs�3�~�K�k�8Gt���q�:��p5�>ݰ�H�\yHk봘�T����)�ȗ��zC��Ĝ{wΥ��;;y�[�{/{a�i�3'E�V����D&7��IKe%���m5]7�� ۏ�A�r ���c�� ��f�?r2��:�U��bJ� �f͂e��	 j(>�T���@giX�h�B~J�|�ABP �? ��zN� ��AJ�!��%&ԞLQEd{Wl���!���})��(�=�$�S���;	7'M�ƴ�*�ޫz��:�t7��TMF��S-0\�$��q����Jp�q�:U^,:�o�:<����(ؠ�����?:�8;"P�=]?�0a�\2��(��|$�!�ѐ1����6��p��������b�����+Ќ=٨�A�	#c��_��$��2Hr����K�V���A!�o?�#��xP��k��������q�$BF�J�4��1�L�M� ��)E�I���푵.h)�%�Ac�cm+��>���+Y;�����R��='6��S��}�lX�b�p���;Z��Ӥ�mMKx4�?d`%�F`���S�:o����O��l1$���C0�d���+���[��������加E��N�?�����?���s|m�:�{�M��Ĩ�-7>�e�OD��=��I�d���"��fO��Hn;F�!��=�v�n뿻x���kC�:%��*:��3��8���� ���ԁ�ۅ�����yT�/�y�=�g`a�@�2��l���%�2�Ȇ�W�%�Y8�U����/@�r,������f)�ȼ	e�P��@m����_�5?�v[��BsQLv@ޙQaw�C�<2��
�C��7�h�?����:��f��G2ź��[�!6��bˤ؊�N�ư�����r�M�x��A25Ƴr� ������;q�X��0��tMk�K��ޟ9`��k�'�E���DR���K�x�~}���ƣ9��O�q�߆�³M[&�0v~�Vz�,���X	�GS�8��|sw�/,�a�Eg���7iv)�m���0Z)���\��mS�!��] 7���_�}�`��; 2x����e�����a MW�W��Ti�j��}��	�3c��ȑx�I�t\1]�u��v��W��#�4�):��B6��������G�hĘ!������j�
�dc@��#��A%�M��"���� ��Q�	�G?����^f:�꽋x���)��[�`Q �C�޴}Ei5��uZ!���34�}���ow���f��z7*Hj~��*Q��s�erA'e��������z�������i4�탪:j}��4bp���ClLU�R��ڀe�.Q a�*��Ѯ�����4����Ι"�w�H��j-y�i��	�''vG�p.x'Ī�36��@��G-b+ :&a���t��2&9�Wf��f�*ӊ��7!c"��J���["u��p�R8��:r�5�#1�hl}O��t��#�&y0���I.�y�k)Q�g$U�l�i�ʡ�^[x��;����nYc��i8��Iy#�X{�F��-6���bω��,��=,���,@�q�$9eA'�u?��!;j�oQ�p��.W\��g�_xf�"\�X�5��즲���G�����X�� ������2~7J䂭�6_��#���L��<q#�jD��L����m��:���N�����C*�������	�[����9��.c^	goVl����fѣ�W4�:�H���]��)7;@��:V�Ѓ�S�ւ��H{����HH
��p~����XSkΈ�|��k�X��s�ݿZ,q����hi� 6�S$_��)��c����u�섮��$@ġu�L]��+�7D��� ����.��h#�x6w�^>����"q�1ut���Ńa�ʍâA�z�Ŏ���a?���_5����	���=�/���`n"#E��!g֢��v���{�	�}���#؝��y{��������U��f�oO\x�5Ѣ���
/?/�Wƽ�`���N�f�M�A��!�b��6����2r����1����:&B$]��%���
��4*Y�p&�|6�+����������7T�$a��}:��A�:�����("�4����s���3Q�z�sz��?�>Ѫ��i��Ĝ�C�l��ޭI�@O |t*#�Ko|�n+��O2��%�߸~Cℋx�N۹���@��^�����ݹ-:X����͙�d(m��i���`P�'l�hװ^�A�}����/͟��Qx�<�y�
�!���H�.��IV�,SI�� �c|���$��M����ɹ_v���[�:Ou�Arǩn{�,�l�K���ݾ!�3���RQ~�#��u����8k�\x��s ��\�˭S�1I�Yi"&��[o�\%�_k�8����]�b�i�+F�Cs�HX(53;��4�Pj�,��axO E�7���NV�2;�op���(?��p�E�����|�+�a�v�������K��@y�F��_Y�1<K����A*dxX!K8���c}'�&ˍ�|F3W2\"㬔ǖH�/�Iѿ���=�Nㅩ���櫠��0�n�B:������;�ܽ�~��H�����r���~j���}$Cc)f_a�ͯ��^��3M��4�	t���a��]eٚvI%e��N�{��z	\���ֳ��q/�a_��0��8w69��S��	
����N�[V�f(W�ri���t�R�W��fc:u����u�N���4�gdQ��*�����Xc̼�%#���9��~�E 4��)�Nb��d���R��k������-Ԛ��D͋�K��1�U��[�$
!�!%�����v�����*���<V�N�z.y��X�j&l~h[����l(�R�D{�vb��/�}�d�La�nm��t��;o�+��h3��q�r�~e@�e�t�t:׃q�L�X��U��Bܖ��T6Ub��I�Uq�����1�Vc�#֏��)�*� ��U`O�[U��`����%�cDq+g&M�'6M�<M��5��T�(�pv<���TX'�"að�	�K���,3\Z�����,c @�O9�H�jt2�|�X��.)_�
�\]��:-�J��k�)�� P�����}T@�%s��k5SaʢlZ��Q���M=�����e�*/z�$fG��gB�  �P�����|�e���H�=��I�\ZXlxVHYEB    4f62     b50�{�X ��� z		��-=)+c�u�K��w�:k�M��bV�����V��:#�</��k����,�8�v$��h�d�>Ċ�3���v#�0 ��ۙ٢�}G�CiI.�)�lL��(kr��-����9$�m���P���4Qd���	O(QY�a/~��h�PL�zy�.�����Y�0ָ~��_X_+P:iY��r{W�KEl���Y\[�n��Tyb�v� \�h�q��}�l�Ьh!}LY��n�#���_�,0�k�^7r7����]TJ�����([��W���@���ۥR���O��\�����G�D�����MD���	r�!jɛ��̠�u;��<�����9���_��Eh��aj���;Ĝ����"0�J��웨2�Z�
��#�@�Ů7R�=N�@�3�����&�cw�!�A+/��$�7��K���4������6�1`�B(|��gZ���˿"e+F�p.�}����E�9u�-�ί�?���N���Bs"a�
:���0���~�)��,�.Sv��hK��r�����mj�U�kGD�9'�;O���aiiu���'��u#?���`Cn�;���Ԡ,7�a��T�0*e����Ҽ��ϐ����m�\qG�)vr�ni^!�L�&^�$VW�	h�~9�i)�19�SK�����)�)3X(^���_�%��+^�-�����i�d"֞k4��D�1�+��,�s2�zJh�q�T(ZU0�U�G-1��t�����A��^c?�>7�L�1�߫/��7���c�v|���'�T��LM�q�8�qod�h�h���T@�[˙�'�ĉ�E�D�D��p��̔0ۮ� P���+A�v �Jl�b��)���L+Z���MV\(�Q'���-�R��V<�b�H��y��m�����#&j� T�L45��g��1����ڢO�L.��������ءqZ�3�j�z�;�A��%SE�;b��y��p|Śf�4pg�ԚW*Z��g��j�t�2���/|m�ҽ���Κ�e� ���۽+=�=Ox�GA�##�뽖�P痛S:�*h��C�2��ޗ�)c���.8��<Ӏ�Ud/-2�,�8��@�n7�{�'�ۃ�T��O����=N�if�Ӝa���BF�N�7A�lE
{�B�U�,0�'I��n����qn���|���w�
@�ٕ��St��[%p3Q;�Gdr{�����Z�¶°��˸��b���O<�����/`4�:ڜ۲�ϋ�]����ѳ���"�J�G���w� ��Ƹ��h:�#�'��,����-^i��͚��w�=����3Mp0�0�d�@��+�|��K#�׸����Nb��Z�<�f��҂�9��f�Uuf�>n�#?�QB_P��Q��qRZ�4�tZx��l�d�S��zE&1�;55�|��#P e�≕{�w�j���[Ƈ���(���:�#x~!I�/��Ed������<�}�zMt��[i";�R��&����vdEe�mr[JE��_���ʜ1���C`�5�q�Lg�����3��>΍èy��+��q�ژ��	��i~m�"TeK27�����O.IN̰*���sk_Z�#9- �:�d��h�N�F�b�hx7�zt�y����U�,X����=O�&d�sV�~��w��/�1�C�_��&E<�P�J�KG�by��]Z/�w'�8�h�Hk�(���}u��I�z���6�
���],�x�k��Ź�O$�'��W;�DA���m��yBS
_"6��'��jk�ik��N��CV���Qi��}r++���M��[�?�aOڈ9@@��O'Q*ɝ��v0Vg�/���AČ��=a�؁�]�M�H\`M��;ItHl��S���GRm���������U 31_�<�7|�[�Z�ð�wh8b�pr�y0)�d/j�熵��]i�X���}��j�������B7&�E�g~ql���ќѶ�$�F�`�>�&��w'��Ů����iZ@b�/�8�̍��ĴV��Қf�
���������[��z�9N���ߙB2#1���F7�LO΂v~6�j��剤�ۯM�Ke��m�����J�m��ۂ��^D�����|���$���5���k�"��(߆;�nl�I&��kR�f�up�i_c
��%��B���G`��l"��2�k�8n�4ݜP�ݺI۝f%�|޸���H*7Ob	��9�xG��=_��]�>#��3��kd��j�kנ���HuU+A��9�|���	�t���0�[�6��]taI��;��J��#�P�u�i�3�q*�]F�z�< P��<��-��|�?�)�\������~Y����	;�5R^���[�X4��Agu�S����ϋLkV��2��Z��S���<����Z�pcH���Hcwq��6��P�@P ��T7/��+��GɆ%��!�F���`�&�W�s�3�!o�v?'īj0	v^yt���7ve�8��y�K���o�&km�~�]�^Ϋ��&K����%����_��v�ϺQ����^t���f��}�Y�);�\=Ǡ��1qxY<B�޸��J��t*'Q�R���9)♉�2j"{5�Ş�t�C�W������ᨏ��&ݞ��mX������U9b/bEc��KY~P�Jv��lk֒Q��r�I6�oQ�Շ\�Y"��$�>���̥����a��Ă��}�}}�7̗� \2V~p�4��p�e��\�hO��Љ\7R'��8�&\c��$Ϊs��LҺ�_p8�Ɗx�9�H���F��?��xnR�y�;q����Y
���h�8��g�B�