XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kJ�X�E�f��u4��_�ϫ��U�8�b
����3⭒�o�I�iD�Uw�P^ǫ[5��� �y�"V�y����v_��z8��u���M��&�A�_���q���Q�=�2&p]�^'C��P��_N1<�����e�����,M����~��b~��HE�Դ���̍��)%�T��7iVXl��FQ��O��ct��i�V�^�C2>k#�GmMJ�7�ȁ4��nm���fA�F�y���[�;rܓ-8��_53+/��~"�>�$�F��ݚ�ř#	���L�^�n�7�n��<c\Z�����Ӿa��S��7UśZ��gM$��Q���n3m��86�tH9��SC���!a�m�;F���0?mX�� ���D+�.v�A�Y�s��k����lIt�O\���<]��6⤇��v+=ө�K�@
�mfs*L�JD|�[Z�oѫ���gR��=OP[���<�Ëݸ�G��t&����JM��o�Q;���s�~�<�}�?zww�ov���ҁ'��,A��K�..�dB�®\���@��[�c���Z0y���]&p�|F��y�&>�>�e3����ç�|D�Te���uHߋ�MH�ܷîa�I�,9��̴�3�,c�	��"} g	b,l�����
e�T�2��E�f��@x�U���"���ژ��U��������	x��#&����<N�R-���9�5��B���D޺0�"����Q%m����D6
ϵ�=ڕ*�i�u��XlxVHYEB    95d3    18d0<=�h����*����Jl9�'���3 ���[$��p���?Mx�F����b6�Y�_+����>7'�^��/�2�i؂�������R��ꞅ�Ic?�0:�#y��n��-^�l�hL>̓5���Cy��|�o��!������bq�E1�{�L$�΄�$_� W)��yՅ"���YԠU4յa�d�����2��_�r���P5���>O�9�vo_ m��x�y/l�Y�����!CtC���fw
�ٽ}�}��,�`/GDx��u�z�$栅Z�ML~�{�pEް�N���s�2�S�膞o���vp�6�5q��)ް�,� .�3K {ʥ-R�:���7Ä��+��Y��^�%a:`� @#���9H�`�Y&B1��[�h�^��mf�Ή�Z�>�����#�g�u|�Uq�؀N̅�k�	���d,.�.�p r���$֗!P(�4!I��_Ӱp��Z%]��ݏ}H���T�s�Rou�=�޾�BĳL)W��WE4ԭ�P9Tꆫ,)�t{��2��F�����݉��¿p:JKW��oWP�M�v�QhI�X��0I�s�8�ܖwe��"���%�:p������ ��6���Pm'�pP	~��b&�W�)�0��������Ώ�$� �w�Y���;W���h��٧�o�����̗Bq��	�c�3�'�w��I�˜�B����M� ��U}E���ŠqȲl��[j#T�@bX�� �}��@{�Z^y2�5����"k"%@2��!g]��H���P��s:ʫ�.{ҡ�P�LU&�-U�f�Ue0��JB4�jt��g�Z8��"�w����UQ��6R4\>�B�S)g�������S�˔�fP�~ay{sT�������ޢ��J	A���� >n]���ʥ��包���_T
7NM�]��������ڢ^��Ա�n��s�Ķ�7jh�����qtZ�I=S23e�O������� ����_佅�EQM7ǚ�7P VR��m��iS<�gY��dkB��">hͱ:lj
��88�9&~��bE�n7�N�����5)=���
�Dt���M��#�Hb�Y��C����]_~�ʑ�����Q����ܭ���e`Rp���f�&c�����[!��s�;�*f5B_7o��I��c�`�~!�bGۀ��!����
pSKR�������g3���+��O�v�W��uix��WWR� Q��s�u��u����D��7B>�Z���ǿ�+�6�r��OT�
���Z{�?J���b'�L�t�|�գ���\�L,ƳS|'0y=_q.M�T5����d�@?1�*]�I1T%G����O�ḻ���=��w��/̝��riS��Z���o�+����.@/��ܡ���Ȇʵ,�yƴ3�FI���A.�\��q�󬒚'���.��rf �,JgPz�y ʶ�k����~@�aYt@[C=	1�����2=��^ƞ�����5Q�2�{w��)S�#�0}h�)$�����C�Ț�Տn�T@����a��y�?��!��@&�9�c63M;viɻхKS�|<���l�\"Ea!�uC��t]��V����ms�`뺶����łԩ�ƛ��4�; d|/yu�3p��#��]�e����.|f�&�]�����A��|#}ۣsM�pX��� �e���˕G`�	�QQv3�2��{j�
�)���cDdQ,mO'�e�l�&�_2rxk\���p�I뼌*�˕{)�Hý�B�B9�\��~X�\����/'��RL���8&��T����2`)g]]bj�
n�ST�hھȃ�$�y6ǉ��R����wR$�v�I<��G�� �i��qB�T7��C|g�sN�eE�F��p�A֜��s��N��6��w����}f�*ET��G�N���>Ȍ�^�!�*Yܧ�s�<��?�2ړǪ-�ڀ˓w�hn��]۩�:���#(����9���I���ᣅc�]���(ة8��ΙVG7�9����;�y���
o@2��	D�?�@-�ֺ=�,]c��&��HG�!b�:��m-�:ʧ9blF�{~wO{�ȑ�s�t�fӣ������!�����J\Uٔ�M���
i�0�hY���]�|�\i�'8�4�C�,�<���ས�A_F�����0'D��,?!^6��C������J��@����ۧw�Sՙ����"hR��8j�C=y\�����a��x���+Ǌ�)ȫ�A��;F�k�L9��	)�X{�"��	���9
v�\)�9�@���襓K�h��)5h�8�Lɴ`�Ɵ��I�N�Kw�����Y6��n�=����;�I뗄�p�	�nb�A��/�#J�Y��|�;���t�z�l�ݟ��Lm}
�Ա�/r+q�T�V�������[���qڄ�(�:�0��oC0��7��E��z�ξ߮�ՒSB8@����0+�� ��F� �|g2��r|�r��y�d�N/�@��X�K2������c� �A)�Q�E�aА�vƾ�+�x�kG��k�eyf�ށn_�g<���܁��o͓�qM$���Bz"7Z-�|�v���pϲH�X���)�.�q����0���ݱf�����\��� �9�&�z7�נV��/Jh�������9���d8���ܞ#38�`��Z1��vh*/{������=>$���"4��_6�$|��9Y�ڿ������A�0���}�����<]Nhl�:�;<>آ����8RJD�����">�X(aL�5)U�7q"PO��3k���1�2����h?�f-�&ȋ���\k��3����s��PݓtݯjA��e����͊rJ�.����M\��Tx���.Z�&ЧzO(M���{k�j4��;ɔ�;�"j�_����î�C��7���ۡz"�� ���x�O�F&	7;D	w#�F���p�����1
������r�e�Ä����v˩.����K#�J}[�j��^um�r��-��e!������؜?�jW7<	A8�='��#����O�c�g���!I�?�!��p.��N����fc�{�pk��1��.�ݦ��^��3�x+��w�����^Ҿ1J ;g�8c���Z�B�R��Y�����o�w'÷"�n'x�1|�Y�`�Q���?�>@�t e�mP�"z���	���ޡq���l3��0t~�?�|oG�U2��x�nX q��uZ��l����HHc�|J���d[@��9d�����,�����m ������=��7
��~`\�!F�^�ħ��q��M��ω[� I������ �-"V+�8�㉣t�Tؐ��;�y�N*h���8�sb��#L^Y�mf�{�0��1+Ej��D8<�o�@x����OV�<6�S������8dA��~�#c�.�?o�D��&eqŴ��{>�c�.�^��
J]�б�y),�u��T�`��߱|Vhfi����n��|�`�-Бrb���q���V�n-�m<SWĦ�`���~݃7P˓����#-��8H&
���j3��7A�Z� ����K�[���~M�*�p���u�l �}��T��P7����.ɭYNP<l��~�8>h���F�R%�6�,���E���oz�·M:m����6zO��,��jM��3S93WK��f2?'l���X^�r�Z�HB̈́���s�r��4��yL�X���_�G���Q����%���/)�A� ���qMf�7}Ӆ�NK��Zͅ6��Bv0�/<`��"�.���S��H;�4��KT�O#=-�ª=lP�.$ߪ5!�PQ
�3�o�V����c�+��W	�rM���~��6z9m�N���t��ZP'��?'(�t֕��_Va7q�w(/��)3�X�撇��@oƖN�3�H�~����e��8�����>��o��,i~
T�EP_l�#�i��h�'�F6M]VUKa�U��.�k,"�b�ew���6_c&�:�H��� \eDr^
��2��\���&��e��n5�XY���0(O�Dw^�<��8n�H�=�M�xM�l�����C�_��.����WR����
fЋP�����V�@�1n?�)Z��t�'-�j oMգ5XF�12B���>�ȭ������\�ow�sYjzQq�&�\��9�iO��f��MY�2�*1���Ǹt�䴨�����;�*>��DΤh,����Ek����S�V�7�Z]�N�h�eG���G�h	{�w�nt9�$�~�&0�qjji�vDIFF���&Z\�"f�h"A���v�s��q��-Q���ڞ�L�/��cLr�dP`!I�$HI�;��	�{�==M@>!n���l^���0^�s���ܖxԸYv[ހX��D�����߶�$K'S��w��vF(�q�ͨ��[�}�[��G�Jj�"{EA���r����N���q?T�w���~�H}����a��c���q�Mq=;AP���?��Q/!���za�w�r��6�-������A�6��,��;c�5���;��̾O4�&�	Հ����y�=���L�;Ԟ����/6�����ޭ4?�J����M�]״,�a"��U�7�����S���0Y9�T[�b��T3�d����f����zG/�NcҊq:��ȴ*pPי����0+��K� =t�k�Y���c1���6*dݨ�U<̇~	�&�`��#ia�"��$���ˡ�2������J�x�Nt��X8V˝@"�?��Iz����ϳ��R|��0�)'�Y�R���Q�"�c3��]|��\O�1����N��U��i>+������S͠4<V32��w�����������~�ٹC=dC߲��F�� ���j��0L�,�#'I!OD+�J�(�'��,�$��c��K��&(m�d+\!���,�1��]���)Le��՝nqu"�r�H���uZ�cӄaŕ\�S�����-Z�����_tԞ�;�	��biX�j��ɥ�KU����M��Fnk��0�c���H"�41�cD���6?0���+��.N�LC,���KS��H��3�7Ȅ^y�t�j�9 ka���Z0�o�����eb�/AwX_�]a�e���ɕ)S�IiV�FY�2�@ᜨ*�2E��'����9e����d��c���1�}}&ٞ;ؿ�*Xf�휍15��4��B�J�U@��F�!Ĵ-~I�Xd,z�צ8�0s�`��M�6�w��Q� ��f��Ԧ���ȅ���I�C� W{���u��c�~�9�xq7A���jsG�
�Ya�T��P�^u���M�#(�&�f"��[Q�vo���@�H�z�$�(�	ijx�j�Q�^**7�f�k���C�ǹ_��hb>:�%$���#1c}���>�6a����^���s�v��G��4��k�Yi'����Ը��1��.��j̀�*K�}��r��z��34�Wgj����^� �]k��0����(\:�H��!��AyqK���Z���5X�ySd�Q��BE~[W��2ǥ��(S3usd)v��0�+kVz��}����d�7�3�_
<-���� �Zl�M�a���@��!��O�F�6	�����i����"�V�*���>r�&�D��W�$���$op ͅ�����~���4�-�_�����w���[�lp��U��.��$��� 7H�����>�B�#Ł�/�єO����'9�
�fmMIf�^B��'g�-�n@Ӥ���|��g�{�� .{��d����X`b]�&�옧%���S�3�c�O48���H�"�9k ���-��s����R��S,��7��i�R��uv���٦0\P�iH1_W1�pI�͚֟_���2f��gi�<?�u�:�dڟeg���Jp8�t6�,T-ʎ�@�Z(�cۛRk�n1��Ǝ7�ae|�~M��T�ev��X�ѳ�Y�p�0?�W�T�&;�ou�,.�$�
J+D��@������3�Ge�v���V��fe�Tт������Q�)�9���}j�2��(�f�M9n����;����7ʥO�?�����?^+��ن�	�[�+��Z��6H��K��C76��ܛ����� ����q��U�eqj·|�.N��є�e���t��c/��O�;H�mv�����(��b��i����߹@�anSV�(�Jm�~��|���Z���o�I��`��o��)�wnzJ�B=%���"�OiPa���p:bi>@=y_�'���7=D