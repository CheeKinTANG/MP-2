XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z~�N��o	j���=�o^K"�	�6���<�T;6)�1G�p�q%����۔7�)o�����g��v*�1#�z{�SbTK����P ��Dg5w܏gM}��Z �s�MJ��$*��-%�Y����j�m ����)ӾhSm���d�䨫*2�S~k~Tmn��w�q:��hAb�y�
Ev�d��U��8tF�_%T'ҪE��?˕��%ȸ,�&OSx.�+f3~�����}�'���'��#Y^���:emr�1�4"vi,9�?D	�D�cq��v;�e09b���)��N� �����^�ΦVw\���Y��(��:RcɞV�2�h]����RM�b�}�|���U��bՌΔj|c߉�v����R>�(hK�RP�D�O�6�y���J�rf��(F��l���y(�p���oZLeI�op6���Mf�6���"���+��'=}-�����0�6��
΂�����ⴁO�/\���^����D��{g�d�����V�V����}3~��~�ֈ/ON���.���8ҏ �r�X���۳��iX���H�%U�,��T�k�����k 4St�`��(�.�R^%��\ZXCx�ɞ���m�J��un�{΂[i�6d`r"��-Eg��b�;�
?�;wp��Q��9�� �c� ve��bS�J`ȒD�ot9�ԝ֯e���C-��?_�M��N��������O����q�.(��)�@�؃�k�|=�T�[���F�A��tGK�i� <=�[AXlxVHYEB    dd8f    21605SE�̸�����8$F+����\Z��'V:g���V����*�z��J�d?��,X#B�1�J���Z@3ަ����]p�_FQ��4pO����m��2�� S�R���H�V�+�
�|�B���dN����F�5�!ԽΊ4��i4��γzWJ�-�2=�fL�<Ҥ7V]6U�9�7q㛂�ت�@PW��;p�5���d��+R>�����S�?ZF9�:�U��_U�aI_���m���p�b]�a�+I��\�u0Q�a�`�V|�$1C�(���^ݗ�˚9��T�fh-ܥ��X���6�o�4-�Ҭi{EU� T�(|�$���Ty~����_�ɽ����m��u��/�P!45�Q<��'A��^��G9�YNQl#����j�N���$PR��]Y@g���J:ʁ��`	?ӈɃ#~�{� ���夠*>�A��l�c���P�i��_�L(A�Ή��;�6�Qc1�	�ʻ"	pEk��v���Mm)TY�{�L�E�z�{3�}��k��MC�������9���Z�b�=�I��{S�Y�ΐ��ӡ�W�[B�@����K�ó�*�H���#g�/�*�>6�npbC���Vmt~�����9�O���Z�8��
��!2�5��B#�i-�;��7��뾄� ��f^S�>=���(m�\��؅<�.@���n35;k�f@*J�
�_�;aG|�'����=Q���*&�����?��1ً*��x��&����ʼ��q�[]�˙v�4g�|�,�t��^����Xż:��M�طg8+y���ȧ@9�-qެk��_�I�1�A���u�%#����eNz��Qm�w���'r��y#��>(s��7I��MX�F���S� ��Klφ�����������?J ���0�#�-�y��`Js3o)�A�E��Y�N���_[&��I5�@Z)
q�62�U�u:6�?�M�w4�a�s��"S\���L%Y#�������t�7�{�To�8�d�WLZ�w�}�
���K^?J,��^�0�����S����|%c,(7x�Z �
�nw���8�����Nr�cQ[g9�xC�/�4@Neq�rn�v�Y����hz��T��X�<A1:�]�܌д)�ez��$���v���s�e�d�������̘3���،t��5���ۄ�������[����hCp��]������f��s�7BŸ2�Ш�o��d�1�eu�K�[켤�'ħ}(�|F!ͩ|(@F�/�~��k�������u�'�����
��H��oWCDL�v6C�R�� [qi�mf9�r\�O�ֺWO�v���Ƙ^S"H��
bb�f��>��ħR�=w�R����5P\ȴ9]��J��o7���|���П���%��T�ǹ�̊�s�����K�/���ЎYX��?�6��U.F�+(˅}
T����&��3u�!Ƥ���j�*�k�3�J"���V]t�����8�<U���u�)�5��"� 1˷T�d�*�X6М�yς�p����ɴ�V.�S��XJ8Rs���DD-����ͥ*
Pn+*r.A�~Ee��E���9X�B7�0h����������HhDR�\�*1��/��'�HY��[�"Z����Ǯ+� I;��0�87@� q�M�ww',P	��/�I-�)���Z"�?�	˳? ��ޟ������IUW_�j�i���L:m������]���.6�4T��9��mV�7q#D���ۂ�C"v�7��6��� ,sEe�ˀ�JR�����x�/ �À$J��{9Ǹ���~%�I��xr4�ˆ�.w�W�� ��Q��ڳ�Z�8O`Ԣ:��H4��h&F�ҁd(���S��Oe��Sa��<Ơ�3?�0ￔ!V���6Jm��� ��}�ɵ���ծ�����.�����b��AII����#��;�x�\�`�q���*F���q{d�.��"�Q�5�/�w�4tT{��/��t��b����������#��ܼ\q�*XYo ��v�<zpm�p�~S��:]���h�u�t�s�:�T��ǃKo�8#&Fo����Lt?�:�#m�q���@~5Pt���k��)b�)ؕ�v��1l�{H��<���=~F��Mp4�h�WoV
9�T��[��:�ze�-(H�B�D]`�Fx&vlX������U݈���A�&N��%��p!/�����bF��H;`����W��x��b�y��R(j������ߌu��杬�˿i�� �Gˆ�e����q�"��ˣ4� ���_�tn��ߟLO������d/ײ1��*-6�p��wU�."�{9���~�=QM�]��4�VfX�F�����R�$�V�d�䋕�:��YΝ6�k6N��ԋ���<5P	"/��C�������E%tL܀���`�������W;T�_��L"�Ɯr���ڗ�/}���,��a���l����>o]���[Ǉ�=��Odwź�#�Ɛ7�s����ҳt�QP�0�Cj}7��:K�:u&�%�tJ��;�zD`p��R��j�5��"�*��e���1M�ќ��o��+�uw
��@�/O�Hv�>����W;���O5��F�y핖U�ZG��N��r\wz�m��6;KYN�wω�2V�PH
��p��J�`ɫ��l��.��� ��8�LT�w�aa��E̔���D��U7� �M�`h�&�|inG�Uu�!f�u����".0�����2�&�u����HY4��b��V~�]�� �VGp��B�@:���� ����yd�����q�=�Mf�W����.ei�k��}�5R�tl"a��o>;��%��o��P�-Pb{~��<w��	�qXj)� n/[��!���˥�;���RZ�.{�Ba07��f̻Ss%䚇����n� j��t��а�p��95=I��4�,=�~��z��P�r�j.�d|��_�n�Z�����@�-J/����
�G�d��-�_���B���������pϨ������wM�}k��xWg��m�WQ����h��k��-��&��uT�{�`wg/�3�� ��#@�q�L(7�{P�䟕L�}FٓQ���XJy�v�w~��/�.A��6���Z�+Z;�g�-�p��~���=^tkv܊�.�����Q)	�q����e.�]Oq�:FA�����b1+\5����ؽ(�V�$ďޣ��M���-��vq�
�Ƙo��^��1��ԓ\�x]�d�q�	R?�<��ʥ�-�� P�����u�g��|�0���I���^�ҭ~�*}�&��>uK�[�PI�:���>yz����Q�S�"l��p~�2:�hĂ�Ӧ(�9����ÁD%�j��h�<r�)H���= ��)?YEѷ�`U!ޞ����vx2���ۭX� �g�&�fւ��4����5F�C������R�g�G������Vȧ���k�w���r���h}mn��p�c�C�QU���+c�����s��ς_Y�>e,_�ȋV�D�E�k�j�4Bx\ǭ�c��΅SY�ȿ����z�o�~ۃ�W��<�>4k��	C�wI��U���[�cӶ#�29��ʩL_�n�B!�k�������a�pFY����S�U�v��ki4ʕ�C�T�j.Z
�����LfQ�\���78��b�,P.�T^�m�ʨw�*ʗ�B��^|�3�cU���T7�8����0��O�GJ�\�ˮ;�g^.�@m�L�G�4��&��=Bw46�!����Y
ޏۮ"�l��9�NO%�s3���Q��P���]9�����
�Դ8��(q#̩�z��랫h{^����f(�_g��g#u��4T*�Ƕ^��C�XyQ1dCS�^�t$C�q8't��4���<�6_Q��LR&�4��$�!�J)˄$�E�
�P��� �v}��-��FS�������N����F����ʠ�3��9{s��N=a�����[LX:���9�L�{?��x��޺��ȽV��5/�S�C}��( ��-9G��Q�bo�`��W��ͯ�U��Ϻ9"ڄ��	V��^��F�"O8�$�J'�ڛm?��?���'@I9��	*���Ll�p���!W`(�:l~D�.`�	���fB*��!�$1Y#�u�!p}G���`�.�OZ?�t�&�[���H��%V=�X.���ĸW,؀�� �!�{�AEf{�2?�q'���V�mB�����$�4�$ԥ�j�c��&�v�>�݋�?p�TvRt��[�@�E�)��4� �ć("t��Z���b���N��������W��������&�� ���Q\c Vʦ�{�iy�-<�ʭ������(,k��.�+;�29�t�N� � OQX��'<����|,A�KGG�P�H'^��� !�Gpz�h���ܫ�m���W��6؆߫�<
|%���A�<������3(��w�.��ke�\���Q�H��ٞ�
��[xC`�=�uZ����8o��
��A�
�a�%8e��-�VmzZ�M�$;z�E*�pu�M5��Z�i%�v��٣gt��Ϡ���Vl����L2�a�!J�hp�w�&����{nv��_��!��
R�^W:�Q�:?�{?j���Z-��V�-_�p2LI��k���Z�5x��m�şB~��>=%ga�H4/JO��_��0�����
�l�(����K����tO/a���(N�V5�^}�$�O�9rt�Lr��?��V@L�R/�б���?�wI}�<��^*�<��Ŷ�h;>�萙KqW�6CP洲��zr�6|�����t�r�U��WaRXĬej�T��	����jZG?��D|uM����Ԩ$@3Zm�مd�ud<l�ns����������y"b�6�cP+T������{xjQ�D&ߥ9�;�*Cٕ"��(@�EcU�j��g���@.ȫ����r�'�N������Z�-��Zs�C���������w�Ĭ��K�gv��o�3�.��b<Gd������nCgp+�Z}"����v�G0w�-�T�*��>i�D�P�]���3�8�l���r�_��>�9/#J��Vr��"�<�Y:|��z���ջ���Z���W���S��1�E1W[`�*�J�F~���pO��ҡT��uf�1_��}�пLq�� x�&@�� ��w���9������J�K[�E(E��A��Z� �uE����)!n�}�&��7��J��vb�<�`��CI�lx����)�7�����	}cc3`�f��|>����}���F�������y���R%�eٰ�xBhcu�R0�T�K�[`'�J6���
�G*)��z�E�Lvn��c�ۼLg|��'zj����u9"I@w�i1�F"�Hb4ΡQSo�w>	��]�P�@L��
�şy8��X�f3�*�&���w;���د��]&��޹N�G_iC%>�e?��X]��I0���z2��E�c��Ҧ�| Q)�sh���g� Mw~=����>�<�J��������;�`�y�wrJ�/'~ �vj�ms�#���	WP<��<�}hv���󈜇<�����\F�ג�H�
J��3U0���U�om����{k�@)� -��Y�d��bZ��vy������Up�=8�W$������]��O���Ԉ��U��s\����P25ۄ����R��*:��;�-:��ډJ�8em�k�>��}��v��U=[�怐.��K��0���)|��{�vp0�o^��?)F{Z������[71ͨ9����I�׵RL Ĳ���j��C�����4ũlTC���va�Gp�=A�Fu��4p�.�2~j��<ьA΀��a�&���j[X��N�.�����Io���sxj��ş����DU�����gUC�	��i��[)?����=�����{�i��$�4)>�:`#�g������R�9��$�֚�D�z41�E�t�r1�w;�c+��o�}�Kի���i#	Z+��.�O���(�i��u�����7����������*�)�*���/�c�-p`|���T���׊�Qu�z��}��f�h3S�S9�*���%��������!����S1�xIe��R���{�����=�#s�eb92�FDl��0
�<+$r��ז\��ɕ��B�����  n(y��������yO�Y��(Hoo<���(`v�.l��a��]��j/��%���y�;�\~M* 76<R�)�u���h��E.�v�(��b*�܇v�C�yP�����M�����w��D��Ϡ�>`|
��C�焴b�c���R:r6��)��!g3� ?���t ����]�R��G�4i���	�����*���y������]�O+LY�&]���<�W�z�(�89�f33Y�s�-{�]5��f��ď&�7��q��n�� s��EJ�a����������}���3���l��G�n�P+]�p��r	�}N�$����tR�-\;�� ��q,0�v�����1$���v��5q�\���������a��U\�o��v����y�A�w
Ă��;��e�� qA��ZZR�^Hb�hg� ��7q*i�sGB�6Ւ{��s.7��ߩT��*�	@�$���p��� F���ٗ�&��˓��x���ٹ/���̫��q�̛ZJ���8�ZM�d%㧓��%]E�7�x�֊���ߨ�	N��Q��4w0eA�so ] j$���6$�FY�G�?3���׻���oX{�!w*�7�b�E�w�E�Uu0D	bxR����q��z��L�3:���|6ا�b��RS�Co￁d�DK�l�L�l��(�ҁŴ_��	`�Go�����6B�xٽ扜�|���6rk~`�Bl�m�L���O��JD"�6��׈�s�I�|yn\�V����)@��bqX��:+��`����y�%Oa��!��7���"��y�
p��."Ƨ��Ip棝������.<d�P�l:ht�1���F��-Dw�X�_���KSե�ꤸԭ�~pB��8��M���ҫ���g��Q���>������~����c�<I�g����V���x�Ͼ:r S��^_0�r]}����ӗMj	��;���>V�QC���hkl���u �g	�^�D��y�3���oT��{�q$��) ���2�e�����~3���큽@숄���A���cW�\��������[M�������T�m�{��6�38<RnɄl��?�y�i)?
}U'��	��CJ�[g<�3���`Z���$«(i���T��F�R�0��QU��Rt��Q�d�����*�YZ��1^rd����qq���z�0�o��5�,�BDo퍙J�4
�ᢆ�uB�Y%˺Xu�K����M�q��K�7�Arl�?/�]�o/(�KD��9��7N>��1�(�*#K�嫢��o sx��:o���M�`��fa��Ƀ�b���s�EC�R��x&�1��wsBfi	#��t������3W&�5ӂ������Xa]��� =�^�r�/�"0��;	U��(��B����h��ty�ڻ&�E�d����T#�4�9�'�3�*�������(#�Qr��>ς/>�C���|N0T圲�E���r��.r�ex�h��x��R^�T�՚Y$Fnao��3&|bk������Έe.��܄!�������8�]��,�{)O�<P�?ь啶����8G�Ɉ��_hFi~Y�5��ai� �XM���Y|�8ǈRD�fy!䷳:��j�E	l+޵�r�#s4����U��UV�]��`=���O����u<#!��5��Io�1����t�r����\.�� ����}�q�����M��`!4mS�Qʚ$m_{��� �]�f���aqF���	`eO�P��I(���S�,& �B�hUGl�r�}b������2,�9���
�����q|VT_�K�� ��cGu��f���S�H5B�-[�	��[�*�ʘ��I=p�7���_��o�m=��,
��h~1e�^��:+(����ڍ�G��Tl6��ko��E�c�8���ޣ�A�J��W~�g��JkY��;�I�����$���x�j����#�Y���W��J�o�b�F��	l�.A
����@/��BU�&��h��%v�Z���G����s8+��T��=N��1қ8���ǳ[B��S����$�8NJX�[$��X�kf�w�wj��������\�;��Y�v�V[�>�@j���,�^��Z〣��F����&�=�ưU��>�*^o�!v��Zu�z��S?����۟y8�m�>��{D�v�ї~�Y���"�Qi([q�"�%��=��p/�c����?�	�N