XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9�nǱ�l�>�#�d-C��}�P���`��.��e2�d�
���mWpFg������@L��I P~�+��ƶw����������m�S�IX�^� ⧣��kQN�Qd}QC��(/Br۰5��Kz�/n�A�h4�`�	HG P a��3���?�S����*uLj�3�p;g���G��;)&���L'��sc�2��`���,��΅�]�I���&hrZq���2������֟�/SXSü�!B �J�\����㐸���8/�h�ר�Z�ϹN\�#X��BZ'/�ĭձ���9/�(���>>���b�b}3���e�Ab�����i�m)��I�z��Q�[H|���K��Ox�8��ٚ�~2deB��t*W����<c׶P�'��i��|ګ &�?�����ԅ���A%�a����0����p���S��o"���T����>�J�L��V7��t��TcVP�pR^�q�%�b���#-X�N�yބ��`���.|k8��G1�~d2���jʮ�A8�$�@<�+�[�6��R�\{x.(�7>��~	r*z$b:Gv*���%TX�"�-���Xj����yU����E!mJ>b�0���J1zOT_�<�l�f�\�����$r�FTA7e�e:��2��[&u��
����H��T�#,�u�6�F�����Q=��g��7mw;�?-8�tn6����a{�����V,���YzF�s���C��%$9�ʃ, #a�_!= �2�s��ɾ���XlxVHYEB    dd8f    2160Sr���tjIQP�r�:�؛#�P�Ԭ �����-�߷�3~��p�.�.]a�2�~A���aXՀ1�FÜ�,-���K�P�ZxRS�M�P�+YO�A[����
�r� ���&����f��&Bxm.�L�͡`�_w�D;�O�������+�%���
�b�+���ruT�rʩa�)���y�u����(��tEr��E?�	���*��@��%�+�'�_4Y�xP�/�9�[�O0���ZB2F��%�b5H��7#�$���_KS�?^;�p�=;l��h�Q�!^���z\��n�8v�BY�����XJ��Q�٩<m(<R��1O��"D� ����>�G��1	&�k�$�VĖ/�ys�nr�vi��<�y�{�A��9�Ɨ,f�%�'����"�����Ͻ�$P��:��`UZ��P��A*3CL̪�SY 5U�m�>�T�	ڼIbK��F����>!`� ����P[\�%�Vd��!e��w���(g�K�O�i����f�)�h5J �8��V��ht^A�rJ��5p(,�g�l���Ē���f�䘤�XN��~>�۷^3�B��69�#k�]�_��+��^�S�f�r�R~� ̏:��G\�>#mї���*�����]'�Q�$��6wͼ�'���x&ǌ �ƊEb�Փ���u�M�-��t��	6��mq����T1�_/�F�$O����ɧ�O!0r�=��{�0���J��`@ER��9�N< �x�k���k"��y�.!2� RD.�߈)���8���iZ�k5�MWQ�O�a�5�Q�0�UtA���ݺ	�X�/��Q_�C������6�V�6�lɜ�2���)�6]�A���B.܌?|��6��0�h�W뺩.��.t�:#�1QS�yb��>d�0^���QtY�iCʦr
���_T�G��˨�{��������Wf��eK�x�z����T@3����;��غ�,�l�:��h�����C:�.��p�w�v'�a��@cW>*�	T���|W�3���'�3��cm�pHD�ux�-@])m� Zz�:�y����	�|ڿ4Ҧ���O�߽�����NGJ4p"�@w�e洔$��#o�^���;���T��al��=�6;�l�
��1�~E��G;�E^�>�SVF�=�]�(�#��j �{��v*[�M���L�R����1��	�O!�|�uߪ;M}����`9)�x��w�cǡi�K�	��X�#;e/g7����A�L�H�+�mPl��m�)����`��y�����I�g����#$����ju"fĉ��z�D�B�5����>Ֆ�@���Opdh-(w6[#6�W̸J��S�@�����@&JR~���U0�ʐO���e�Յ�N�������T�S-v�thT.���>��3�P�j������'�{��E�h��[K��B8+�{X��:�E�s*" rb5����D*gs���V�Hc0���s���L�����P�l�ޠ�?s�o u�wK�~󢮕^�r��L�������s0��D���'�Vlt+�5��4���_(Iq&7���'ľ�$���k�CX��R�U��y[R���M�F?m� ��w{�Z�-u�p�m�\<>�ڻ&i)1��fUN7H%!���|�@�v*�0[�#؜���>���e }���k<�-^�p˔��=��[g&�[S��YJ�Ce�\����XZX�K�Y-���j[H��zI�AĹ�;����T|��Ța/7R'��PZy�_�D]��X^j`���G�<N�~��\��#ѡ�[{��ϗb��C:ti���}U�>�Rx^���iT��(�ۻq,��I�c	 ^�h�:|U�}Xvh�-�ykO�uPEc($���4Oxs�-�������c�҄�x�duM��
v?�d��]�TQ�4I1�h[�m�����F"��J&��Q��	���	���A�qM�L$!�9�|)��@��)p��*���(5�`}�<0��
�'�<~2�S뺰<�j����[�p�����vD �z��eΆ�8ja5�I�FC�i�H�lթa�Q��
��V�Y}?O񷶫#g+���zڸ��]l������i~z/!J���qk���e6o�C��R�1f�9��.\���T���8�?L@Ux�8�fqAwFW��{���^b��<����s!S<K$��H�K >OU��#�ݬpiA�>����>���Ű<�j5�O-_D#�9F7 g��KƂ裐ʌ��ôd ���p��e�Î~�h��>+��X�0EL���A�)�NB\���-�E���h1�3����9W-�[�\?L���\;�jը�I�x��H䟑T�����_�5��W�Vs�(񔘶Ge�v�{6x�20H!V�s%�l9�sU�p*�����E����M���Ww������e=mÉ�co��}:�-Ӗ�ʛ?�Y��x���a4�ok"�QK"���F����ŌS��� b�*,�di&TWBT�`}vU�ѹ���������熭h^����V.S��/�\�s��g�k�����Ki*s-���;���j�̀A�/����r3�er���i|gb��7�\t��>�ɲY�0ʌ��o��ć�g�t���%�#O��W�"2m�夺�ш�~��e�ĺ-��ݛZ�2���o�0C�'.V�9r?��[�Q�@��"TV�j9N�	��_PqA|����Se"����[������c����&���:M��kcT��R�_�aqX�\��)}.�	LH
�]�WeD�-Ɔ��<�
1�	F�-0t�:G-��0:��LV�:e� ��]�/�:���C�a��ω�ңP��N
�pu$��-&�bv�ueܼ��sU�u��U.���X�����?Ub(\��F~��h�nV-���=.����6��ҭ4�.��z�Ɏ��V5�e�U@�����BW����p9�0׬W��i#���OV�	\'lܓ��K�q
Ջ�D&`ϊ���_h�@��<��C�xR�!�0aa��q��Q}�,��]��	��ՠd��4]P��u�\9l���Ƒ���5��v���!�q�n�n[4� -T�\�d��_??5-k YB�5��"���&5��VpYd���N1	��_|����s��i�n u^J2Λ� -5[���@�>�e|9�^������k���=�����/��=ZE�m��E5i�.HX�G�w9I
6�9#�@ڮ��HLG6��*b ����TX�F�����$F��{�~Lp���3�J8��;��8�a��?o��9���$�ޘ��&{��rD-��I*�� ��H	���4��U�c��Kg�1��2�U���m+�3hP3|����2�U�R��0BHrl�XcVV�K`��ɛu��D� ѽ+��"�{Oa��Nة�{�|!y�z��"�ZE+6(.�>�1��EV%�Z�<rߢH8�=XR�ڄ�]!�E�[��c[�P�ޟ��V cV�3���X�瘂�y�{$D�=\]\���<�Ќ?��uJ�_�	:����h�q���Td��u����Z<0��}S<��F�	t��c�37�L��d��Ⱦ�6����Zi��x+DLSko����х�(�^%����9S;�Kt��N1����Qɺ�_�Ѧ�j^P�ȩ.��;ۇ�π7������9��~ї"55�*�i4�V'"��Ri{�����L ��y�1�����[�Oİ�����)��ܟq�?tU �s� ��G��oͻ���@�!�P�z�t��C����
#0ݿ�u�p�~t�UuVOcS��ʼJ�a�q�Os��O��Z.J�(�����!�Ȥ9
�?f�xӏ6f, L��Y���8cjQH�8���n��I��扬��jY<�Ǭ�_4�k�iv��e�me�wE�ϔ#�N�\/�1�f^�5	�JG�A96����>RJ�x��n��t�<'z�mf��Y'�xe�fױ���v����Wi{�8�@����P�|�����r���8\��'�E���}�Pm��E�0�D6,��.�Z�o F6�}�h�~ �hH �I]�%-���K��k��t��Є�"�%����ݻ����D
��H��r�!��P}��u����L�<�&�� o�%�LO/�FI	) �q
�Ӎ�|�|���@��{&$ږ�"[$V�(�Q�|��Xz{�!�?Leyk��z6���	��2ğ�fs�� 7�~p�ף�-�:S��87?y��F��kKܩ�ޚ��nq �A"zp�x!�
E��JaC�/�B��(p�;�����)喝��_!�#f���1���iH�
WVi�?��}M1����	��)���p��θ�᪋���~�]�Cyn�BU�^E�3�z�.����*�8ۙ_�cK5?��:��,_Ðw�#.;�X����\`I���Y�blS�����m@�tD�(H�Jr��"�_jDTŒ�.�VRe�(��'��l>���0������~�(98&w�dF��"���G׮�>������6�2���z��z��R`/�6j]��S�6��\���[Ĝ�==8pxO��7������
h 񂵄�춂�#��-%F��͕������-�p��t[O�[����id�Қ�̎��4�S��-�PgWL���}oR��(L����?2�V���(��M�`�7�%q�����4ѳA�[�$�g��;N�_�{��6�m;��i�`U��qp:��%ӣYq�s�&گ�[��q�r:
n��M.0�kf|i��5?8��Y������[;��i�!�?�������S�N�|w�eF��l��G�*�ɷE�_��Īm�z2�
�e+�ڽ�w�}�t9=$}�����[[7y]VK��t9�V��,���,CͩIGWȬ��89�M]\�ʽ2:�/ȸ��F9F�l��~_r(�	�.����ņ�P�'=���u�P��|��&�'0�涼\���X�+�ʜ�mPH�nŌc\䴒�_y;����Fr{��K�<�@���&2�?yQ��Y��ZuM�)��:���R�uk��/39P)-O�w4�������+�� x"ROhWD�f�Q��Ξ��/��s�h*��� � <	�����4���o�̮f�N%�1��p�(�+M|�.:�9�t���6"���6$��[\��?�û�����^h�Wd�0�������3�o�tF�W3PP�=�m1Bg�Wk7���ޓ�6p�(��u�W�tزK���n~r��/W���Q-	�����ǂ6�Z�|N?<<��}��m�C*f�)E��cDҐ�~�b���i���l�Vؓ����ط��'��<�܎��E3`w{t���2٘�ࡰ�&.W�@ �&�0���f��x��ş�4{��?�
0e"�-��a��G��x�V��(����j��>�m��zj�yp�¿�4�7�)O�TaT 2���;��*����qsŌ�4+�t��G�呖ěݦF��zw��PV�~���Ơ.ہ��E3U �<���К��6c���"l�ղ�S������kHl���0o��bDH�����Iq>c2�K�e/,�*��������i�\c�ǂ��\��G:i�'t�)�KO�~+-E���TI�q쾭غնDy�[�Ln�.�c$�s��J]U�ùS��*�l��,�kJ��m��jD�_Y�"��;���E�苛X�$O�����)�a[�������= �N�ǎz��,<K<ٝ��m3:��X� ����b��k������^.�y� ?�f�� ^X<� ,"u�=�֏xI:0�c�/���"��sgH�~�R�H�]�/�vb4ȡm�p�
�r,$�r:~RG�����a�;d����tK���tY�h����gL�>?l��t,���b�������r����Ikܺ^ߏ�>xV��[�,��&�r,���)��1c�O�˵wP�Y�Зn�y���4�q�Q�ӛ�'R*��LT~O�{�r�i�<!G���x#�6�q��Z�X�R�u��yh��1�ӺT9��Xj���A��I%Z#��D�.���+�`�
t�����8�b��U��ر�Art�q��k�y"0�������3��{2'�U���)�0�(N���\}��S���Sbv�pK�wWn�+襨�ՠ|R!�tZ}L� e�B7�����X�b��m���e�2���<�N}�m�b�ꠡ�Q�oɶ��V��[�N0i�<����
�`��ݮ�K�8�2Z艬��fn�i�D0|�H2t�̈́�����'ޱmfa�ʯ"z��f[���H�j�ep��Ą��=�%��sʊ|��#��.����,b��岱	�<o%�$Ed[j�����&g��)���X���U�$�m�
�����kq-o�����Q,l ʱF�fƱܑ��ؑ?�Z�R�h6�y�����K2�
j=^'��U/�ev�����)Xm�V˧?xc6а'Ig�E` Zw���
���{��=z�r�Ӿ���B�e����ƴh;4�=�O��}�����/\۽��EwaXm>b9W-���w�ҁ<���F����IZ�C����>u��};��G��U���Xi�1���4i��	��^Ǣ�B�-��&5�&v�G�V��������4yvB֣uƊXlZQ}~!�e�fu�L�Y7,$��<`�m�N۽0^Y�@3��8�X&[�qL�p��2\�k9W�Au��2w�t��Ə���/�\Y�N��Rq���S{�Ӟ@m��,E�J/�	u��G�@Hd/e<+g�ItH��܎�y~N.��\b��S�c�{j϶��\���l�k]%ꀻTyۿ��­�M�H{�vf$kZ@�:�/�N�Z'�$�izM�(�� ��amg��]�P���� H��!UE�������완���%�"E�G��K|6��A��ԟ�z�+/L8��&i�u�`�JO>�18#��lȽ8_L~��nq����#x�Y�\v�3�:Ƶ�+��CӨy�I��2����2/~�M����@�o�ݭz:�=g�>�T���l�Q)_��W�����E����1_9Yj�2UE�(	�%�Џ�g�XV��q�b�JѪ_��n���cU��7�F�IM�Dد>e�M���g�S�tH��k�I\o��v��ȁ2v"Ao������D��X���?�.��S�ny��~�#�߸ub���Ek�{�jQK�u�o�Hl��r�~��5;E��Tg���׽�;h7�.}�1�E�޿���^.�;��Da�y��lKY`X�u��N��$W�Ͱ���C�M檊T�c���è�7�~�����_&�Ǝ1rL�'!c�f4v���6)�{�9-2���>'�[�I�����nf
� �
��i�Jj��J�>m#}�Nwl��ӿ��G�QO�:�<��c���c�ZmA3eDƭ��l��~7_�<�T�S��)w���0(b}R��N�����qv�1�@����X�T��)WP�tK*+���i�h4ߘ��mF��e��0�ۏ���~d��X"���Cߛ��t�j��O��$?�m�3�#״O��^���hH�Uv%%#�����A���T����U�Q��7�F���8�g)*��4{��S]u(�D)3��={b��b��N.�߮�q�?�!���3`'�]���<B��b�o�jX_M���'r���/�RD�����X��� ,�w0@���0)�v��V|��a��ok@E �OgN޶5~�Au?���ǅ��}��%#t�f�%���o�6�hlݰ�@\�����M���V4���Cr_ P�-A������j�7���n���o��x��Z��js�v;���B�P�cO�-�,aI�?�a����kM�Fq��O�DZ�ip����~n��,�
p�� e������d�g&�.uSx��ĲOq��.���O��u'Gg&�a|�
�Ǹ\pW }��_y�E�:�ܑ����E/�C�^c�:�Z���13��|���C	�s���Sn�KN��M��B�#� ~s`w6�G���i,�I]{q�q���@�(� 1I�i¿��~�b�ͦᯊ�|�T��,y���o=�2�H?�O�ǘt��z��_ 64��̫ЙN��!f�6�u�F�
���h��~�w9':Į����������?�褦łdi��/�����%2z  �[����	+������-|�BR�[��	_ <��<��ի�lڑH��9Z\ #��$2�HnN�h�	�������Ԏ������u���ZfsA������뀴o�-����
��0�w������c�!y>�?F����`N���32�����R��I�.X�:ud�_�d�6��:�u��=��k���]�����Y����]�mR_�y,��n
yM��