XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>{�l���QϏ�U �,'�%���韧�bGh��ZDj�@�"Z��}���(zceƗ�'s��F�����9`��P�w4�P�I`� UGG�d���M�
WQ�k<�����Κ�]}Rt��Q��c� ��0��k���+�I�Lz�Q��'ץ�W�����=��5���1+XR�R�^�[F��%�/tˆ[?5�$Xv��ľ�n!����,�U���/L���70�T�
�ޮ��*����q*�m�J�@w���ڿ��T݅�J��v��#����C=��<,F��/M�=��/wb <؎"6M%_B�g�#�MB1@�kT�@��W`m/ �=��� �k�T1�������[]c��,��>@k'L�P�M��Td��U{�f4+��k�k(�F^�v�j�MIL�7����P��Vv��DW?f�i2���"�{�F
�=��b�]R���3͞�;�+J�d���\J�H/χZ{�Ȝ�&�ӛ�Q*fNX���,��N<�[�|���r�eJ���V�.럠���.� 4:�D�(���[!����99���ߵ�j�{Z4���\��3��i��
ڗAȩ�H���Fu4��S']�+�;�Ir���1��Kx_wν�������
�6=��������W����Pc�� G�mg��W�rbJ�:��XG~!��_]�t�8��hl����E��@�CQ��r��iv��2#�#_����F���P��N#���Pt}�;�XlxVHYEB    6315    1790��&n���|��&��%���j8�I����PB&�+�Y���������9���X���W��J\՝�����(d�ܳ� l� )z
������'�'A�[?�m�>�)eK!�O���q7*�jr�ǴF1r��!\C��rA����3�E��-�}!�[Ii���:1Ao�\�1(CBK(ְ��]��#�h���N�y���BA���˷�Խ!X5���4b�"�L�)���J8�'/���bi�h��$���tWCQp�g����E���E�����z����b��U�ηV^X+.�����
�M)�2.�����w:�5SCN�ƲErC!����7n��M�s:�p>b���'�g�Ol�2 �K.w��#mFux���)���Ci����HB�(��pB+�B�/~�.�Z��@L����þP#��+s�C��eVW��4Yߓ΁�
����>YJ��%ԙZ�	7�W��r>�:������[�Ϛ�"P���9V�l�±���Wy�U��C�3#���K���=�����r1e�`���#ͅ��^�3��Q�-f��g�m��D>H�գ=#y�_�^�Z���~�(��e����Lt��m2����pa��ID�/�z����/U���g�rp�p���S׶��2� F�v�ŀ{L
�Y��*&�I /� ��a��@�j�<��G�*��?��H2�Mg�Rw��ڬ"k��ҨlC�W��mtA�L�ܳ�@����zf��]���8���)޲<B:  I�d~N��[��#�D���c�Mv ���搔U
�4*��v��'X�%���]��l��՝�����!�h��9����y�)��ˏ�*+Q��u��,n�x4os��\*����"S^&�ͼ��b�")�Bd�~u]��z+>�����v��4\h�����s&���<��x���Q��.\浖i}_!���3�W�&z���N�K-�C����&u��
�Ι=s{{C�Q�[5PZ��ݡ�٘�� Nq��t{Dϰ��*��n#*�7}��=�����`�K�ۈ�*��K��C����Z��s�=v�t�B���R�I=��]*�iXɦ�N@�'̥?��k��u�����[��mR�}=��pά�N~H���F�o�z*2pi�����qM�q�t:�q��k��ߣw�c�5�	��q�n~B�I����b������k�����臿�5�%b��|j|����y������N�~n�ײ���ޫ��a%$���UiEt��\)�����f��V�_=���^�6	��#M�۱�Ƕ¯���L�������=G8������N��~5?�w�C��F�X�Ď�Z���^��e@��	��R��N�ByR���i�;L�+-!��r��n���}/2�x�Bg ���Β['V��']?�'�&���Mn=�=k��Â9����f xy�p����<L�W2c��j���
5�$5}����\�m�')MOɿi���L:z�vK����Y��L4���N a�Gm��T^0|A�D�7�d@����ǐ��;����m�07Q�R���A�
�(+�b m�]j��k�b���FV���0L������f�Ի�X- ":��j��:�z���z?wLE|h�_����Y��.�oY��D�ɜ�]D��`[��}eKKE���/fOV�����`�pR�A��A�ѕ�)�v���w)ŏ�;�T����U��ڀ���~sG��������$������;���@��LL)�dUtL| !��6�2���N�n�I"����| T��'yQ��"%^��^	7d�Ȓʹ�S��	m^�g�t����ʉ��ծK��T��� bd�I,��yҀ��޷�D�'��֠��u��cEUPUiv��).�V���b���p|-'`�/�GgD�X���Jm	�yK3�+�kL0���x#�zB]������C�o}�׿		+��P2#�9�;{^�u�\;-J.rC����0�t���Uq;Ϯ�{l&B�b�2yh�V�_�0%�s~,��+�2����ŧ��
�)��-
�2\���K���`�t `W�)�Z�0;��K����ZO9�ש�4+�h���0a�2����g����X�\�E|H���b,���~Y� &�^Sf��PE-��'�Z�5�t��8W�kf!Z���#�G`��$��0VC8�@�"8�N-_�rD(�%�'�ܲO�%�r��l�NE٥#b���k.�
��a+�~�w��#>�ٖ�A��#eA �~!�U�Dj�\�!c��ļa��o��#T�L��E�ǗR�N
��?�#��Ѿ����UZ�(?�/�R�m	6�8Q�M��J���'��
i��O��v�8lI����fx:BUA"ŨȌ�h���{	iR�}����:h��_Rx/���i��,��y�����Q�ʕN�_�}<b8��x�XPC��*^����E�`�[�V.���#��^U�/�hy#���y���Ԏ�������[e?^��Ӓˉ�\�K�����@|���o�;	�GS����t�]U��k�#�(�Q�?,`
{�5Fr`F7;��pa�t�E���+�KCe��Ĭ��>�������l=p�El�R3=.�����}�zJ����S9
3\h�12�%��I	��~�"���Ke;��{�o����N$ж�����@V����JQ�G�y7������r6������rf|���Т]%l�4������H�ˣ���w�&��۫�Eg*��S���d>��r��uE����� >d��)�@��w+�&/���9��~��_�X��%������ )�p���?;[���h��R>�N���4!��P?�!K^a߹847�\�,�ŋ^Y9��R�PLn�p.�A:9��BE�����m�5}���u;t����c��Z(�vU����*vY�]�e���N���;�H����"�m�v΀�˱�ȷ��a(�E=W��N����࿓5�6ZMjj�ճ����q7Tgn���-2dD�����a'�������	��jO'e�17����)��ˆ7�e.�y��WQ68�R�N��;�K"�Q�oHym��:����\3����֖��>��V��`�&k���Q;q-���]�ށ;b?K7E\aY��{$&�jȨ�/w�+@W���%N=^���z�+��D�-�Y~�3�&|ދ�ΧC!ht�k�R���]��Q���kܦye���2o���~��]!��+���jJ�σx�szMg��t�Kؓ�PS�_
]���tu5{�'�����PҀ��[c���l�
�_CfJ�N�`w�`���v�.ډ�O`#�-��|ӝ��<o疪 ��I`�tAo|�INC2l<�]���:� �I9����o�(tw��������=!H��e"��3 2!M�&.��KvV9����tt��`d!��N������9�Dӈf���/{��̄��u^eF�+���
F�Bp7c����h���ɲ���\Y�.-��z��kV�br8o��Wrx�x�� �{�L#S[�Zx��1VwɨlS�L�S>j&�w�YI��'��~k�!�1*�����̢4�W�
�A�D����nr�]C���B��"�><���^U��(DS`����s���wӑIh�������R" ԭ���@"k��ws��"'����z��>o����/���T�3�����/P2,����[%� Q�,��.���7���B �r,$�P2)e�8��{�|���Z�uJ�s�v�P�H�����;{�@ыа�48�䦸�!���^s�@�M�O�9y<#���+ Ҁ�S������
'x8	� D�.��Z����Ѧ���Iܯ��s���2�>���4P�W�Zva����-�tq�:�iF��A? ��W�ځU_�*uk�ޏ6\��A���hQ9�~SFuy��RĘߛ�����|k�kiQ[H�]ߨ��U}���N,����<��bL\
Pa=#��Hh�e5������kL�Q�q� $�2!�@���&���3
�q^�������`�+�6�7ei�n�C�qK���Yڋ�8�P�z`�M��-��i:��Q��n��"C=�J,�N��:k��<�M�μPUM����B��4#$����~�fO4�U�|�e��3����W|2-�e�˫(bj{ �.|�v!��${#	ui��_͙g�RW�qШ:�{�uڕV7�����H���[^|��kt5�I[�C�8#uLA����Ǒ!���D8�j�#᫩�YDUzPي�ǰ����.j{e�*/uܧ���=U#Rp��B�N���>(��G֎pN/����o}�h�#�K��N	���P~�A�z��a[�,8b��!�7}B?�2�R2;�͢ǜ�Ǩ���.�^�D�p������;��4/��(�l�R�(�*x��P���ˤ��)�QI���H�Of��[YX��j��'Z���;���o���J�pnk�OFe����l�	�t���1�����0c~�dO��_�>�O�y.��$y��Vc�㠵�b���.0��j_]ƺ����Y`� ��wMm_e���kf�%�Ӓ8�[��%�r:��O�JDj��à.[� ��[�qW�4�1R4R�J�Ĳ�Z���9��>��0�FD*Sn���2�#P'B����V!�
<������NuX�w�k`���9UO��7�7m透���'��y�ۻg^E+�޲��^E4���x�"<"�v���w�=yx_ɥ#!C�$S|�	�z�����]�}8I�wܼI����P���j�m�j�ت�6�p��ɇU�8kǽ���+���-�I;2F��5n��*�s��I��M
���З������$7���S�rnt!�˙�i��Z�K������5���9͏@%S4�A66���݄,��Y�.��Eƀ2$�K	��9�t��7oeA
��@�R%�/K=��.�C#|�,�(g9���*�P�Ι���=v!f�ô�N��
� <ZV�*��q�jI����X�1����\bM5��~�0m���:�V��2v'�F�k��L��$����fG׋˂���vSP�����y����-@���A�SVW��d}���#�����J���7�U6y�F]+�oޭ��=	b)6�VK7�]�p�ӡճ�,�@�K��>���e��\��8��'I<Sv�#]p�Z���n-��TbTŇe�%N6ο.��Hg}�f/�D��B�����"r1�'�ͯ�#��,u���P�����9�T�e����6�h��5:>���?��6��5 �h��`0;�H��l��9肘YLUv�5Ruh���>j���x�1K�Vڴ�`o���a}v��"��������0$��ҥ���g�njAӘ����F4">(��L�!ww��{�;z���G��� �G��=l�O%`��Ѥ�� �]����@TB�Y��}�H�>�{��\]"�cNK:Z#/O���o��m�B�\xT�ό-Z\pJ�F�t1���}k�0�a�B`�G��7��="�*a#C4`i#�{0�sEd;�a���h.M�۳Y{�Ѻ6囈��ͥ9��7��5f�_≡�`�A�ͨ�.1�qG�i��;{*e=O`���W�R��+�f� �c2)s��ր2m�-8��B%G�:фL�7����LS�)tI���E���i�u�o��6d_.A��d����/�Ʀ�.\U�R)������x�q�AV$�/j�bP.4gR�Zp?��'�`?;��6{{��	������̨e���ƚo�>�?411U�(��9�6�dJ�� ��!l�,�u>>&�Yk��rƴ���Ru���C̷�Q��2���-�5��[��<L-