XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i1~�'|�1�kԀt���m<޽�e�i���8�^�It�-�o#��AQ�YBv��mF�m0jnXq�\p����CF�+�
M�/����l�3�2%.�?�[����Α�NQL;�&1����d�nfM���%�D���	i9T���4Uu�IX��M��u�羟�k��� ���R�=���s����&=���"C8�"(iE1J�'e�g�j�x �:`����%��s�p	x�� ��d3G(L�b���Q��N7�D�'�z�Ԁ��%_/l!-`{�jd)����#�8�F3��3�i��>aǙ�~�r�]I��5�((PgK��jn4:+��ڝ��H'�L
�s�7R������s���q���Z0)D.�ܻ��sF�et5s�vm<0���	L`y���b�j|[$���5�~\�ԙojs2,��}�&lf�ij�t��K'��e㛳���|d�9���
��O�� Ad�_�MѪ���Z���HU}��g��y�x�k�2�o�O+��#�B��!�V���,WGx�`�9Zwey��m�r���,}N	Jٷw�&u_<K% ��o����*�`��α>�F"�*�q@����3ybMk�l*��6�kLSU���o�	Q@���T=�\���7,�UR�3����mP9��|��6��O�nd�k�ڵ1����jl�2h!��>��&������U��P��ӫ�U��x�p|Tmvav�[�p"�� �Q��o�_������a!m�XlxVHYEB    9fc7    1fd0�Zs�I����J3lƝ�'��[� �0��x�-��)3&& 68���8�ǆ�>|g#���i���rU�P�0ŚU�\/��d��Cc8��"�����dP `k3�ܿ��$&�q�dt%rm{�K>�	&T̛z�B�����w�u:9���!�Bȥ�$��~�^K���|'1-\{��6݊�y*��u'��I�8�N�^@h�r�'À�!�+��hr7rD�	 r��
s<�E��l�|�i��	�]�����j"��[�����_4PD�l�5wɥ8�Hn�P�l���.��TQ�*�mW�Xq�A�ؿ��>�2��uf���(�6�y=���O@�B"�=�؃:�V(�?�T:���_�J��ۃ�.���S6��:L}ٹ�j�}���L{�"BB�)�#�;�Q;�r	C鎾U�1QۻH�@D�^�	� A�������� g0���h޽ Q�'�%�����S�$���;�^9m�߉��qM�����,�[�P�C7'K�W<��#3_�?+<۶$GD7�i#̚L��﾿�f�%�3�`'��v���yZ��&�@p�� �3猩@�Eڝ�5ή��/��^3&ךz�����r��]�y�Ɂ��i��6*.ԡ=*K*$�3��I��E��2JNg��'M���W�3�Ch�oa�u�-ݠd�à�g�(���+��9:��W������b�$�#��>anI6��ee�e 5����C���yC��[L�d�s�`["2�(�c�#�b�~A��A8O�r��?S�GY��R�7���K�����T�a1���첶����&�3�|������O�[���ꙧ;f�2Խ;��f�49�-9�@����D`����T�]]V���]�y�s/��kڮ\��G��`���m9�%�b}㫝�hO�Q��b'�Z��AS"� �/��)x��V���fC�J� ����kS�"���,x<pvC�p(��d�d��ӿ�U�Q~L��i�wG��I�T_Mל
���h��͛���OX�^��&�\��?��7�)J{S h��q�D���_k�����C 8t�,H���u�����_���-�ω���@��
{܆�"�r������������	(�(�ҳ㥙18�x��6Y�$�o�>B�J�30�TX��H�Xrߦ�P���w�ې�����Y.&n*�,�S��H���������lUӖ~���

�k/=LE�����(]&F��db୭��)G��K�1���a]�v����"��<��)��DK�:�w% ���r q9X�����teԿr�Z3X��D�Sx����(�&j�Y���9��J�4U|F�����f�@Q�pk3�%ee,H��z�(*K�%%����myL�`���h�Կ�>z��TO�?���O�׭��ɡ��A�U+	lQ�� \k�,�n������Q�̓n��r��HV�CR���9���͙bdlw��I�/.La���4��� 쏙?�����C�6֪vh��0_�}�.�zE�kQ�ɂ}1�傩���ֆ���Kv��y+�n����)��pW�V�:��t`��D������im�T���Ԇ5B�,�~я�i��`��y)�tB�s~�S��go �1�fI״'�c�S'e�}K����l���}2l�����B`�#�FE��ȁ)��%���+����W��9`N�Ć(:B�T(cr�>���p����n��4i3?@3�=(WuF��jW����|�Ag�Wv��\�_H�:~��J7�i��F7�B"T0I<<)��z$4d�b��H6��e\9ʿ��Ea_4�rDP1F�w��L��M��ޜCQQ�M�&����������Z���ag��L��V��NЧ���3LR��;MFR��?,�������/����B��ĭP��\}�?¸n{�b~+�g@Ӆ���!YQػ6�]���2K�DjU^�&��w�M�|��iɴG��A�!ó����0Š5J*yQ}o{M�߰Yx� ��w���2��h�����s��E�7I�ZUM.�䮰���e=�Nщ��<`�^s���e����X����x/��)=VZ_�%8B��P�)C�&��[Mc�A]��v�C�f���
��A?p��0���&��9�[��L��}��?	���۷���Ϋ�a~�,4u3c�!��G��YDuc�
�C��G��� 뺸�w�<��l��7%�&r�%2�$���因{�7_�%s&��j3dI�Y�X��4�g_y�bJ�y-��.��)����r>�7,p4����Z����oе�[A�����_�|9ƁK��������kj����2qȒ���:�h�zJ&ɡV,��iҷ�u �4����R"�ͻ	�b��"!�����	: !�� �]��(:v�z��t��sl#�����7�"
��G�z��B�M�=�����@��QÀީ��ӂ���q@�ú����}�)��(e����#�Ns��c[@ИV���M!D}1f�>�u�q*&,�7׈�/�Fb�-Vh�7K�	9d�i�_D��r]�_�	隦�� ��˩�_+�.�P�̹F�*��U�ݼ�f<��:��<��k�ޠ�']p��3�Fz�wc%���@��,� T2��%�? ����.�@�[X�*V����+�uw��Y��<n	�;x�>�^=o�2),�	��2���.��{�\ҵX	��n.�j%$�p��LR���Q-�Ƀݓ���b5��A��Bisdo9.�y�\����ؔ{o��Yo��ݩ\l��p�ǟhj�X^�ψ�Q%�߲"\M��7�(����ݵ��
J����OZ���Mk�q;��6YS��)�x�"�xj8�ܢ"��aQ=e�l�g�YB�5oL�E.�>ka0���6���*Q�<����p�.?0�鞩���$�߭�����T�Ҥ��f�����ec?%y����[� ���@�4��B��:��P��8�OF�^& #b( `*��'��P�0�C/�b�����sQ����k$@���p��|#��q����6e��$���gxע�X�TY'�i���`^� r�h�Y��Ы^ n�Z��/��
����m
�`����:K-^ԅ�6S����s��^�;�
D�&v%��~�Ͳ;�,K�u*ж�\$ѹ,�BCR&�̟sv��Y�9��!�'3�;��iB\J3M|r��)��8�Vx��	��D뻇{5S�����`�/h��P5��r]船yn66�Y�[��i`x��1n���TF{b�2���J2�	V*�.�;Xs"���X��W�o�-�i�Ei�s����gK$䗮�`濏u���0P8�
�)��AF�$������5{��*��ک�0,-�Y�2�x6���9o|��G�}xy݌�b��߶'�~g{�OPw?>IN|㋌��rK逩{�(�6�^��eѼ�Ƀ~<Ġ�P2B��^51!�2�v ���#	eOG�cg܇T�K�W�m��d+�D��?M�����[e�ƨ�oʿ��9!fE�<:J��f>���#"��5���!����h��.�Q������{�SX\^�s�(�=�������-�~t����P2��r�+tLn��Q�CXf���r�\�6QqKD�~�����%���M��h[NR`zp���)�虬q3d<{�n�f���lDh(F�������ٻ�N����s7��*�&�Hl���)��j���wmD��A"�nE���Yn\t1*Z|���2F�1h}{s ��u��j�o I�5*��v� zf�G��F���V��X�����D&�ˏX�9p^x���4�1�и�(Ê�]�b��C[�i���X+�e� h0�UKY}�0yҀB�c��-Zw�U	
�����-�zu\�����Nj�Ml-�u����d�����Z&�QF��F���Ŭ]��� �9�`Ŕ��Y\�Aí�-s��'
�-�����R�Z�&���#"|��YC��	��dM�M�"��j�K�;��ݗ�<��ϕ�z��{#��W�l�?k�(�����t �2�%����!S4o�WΎ�.7�"���M�W�˰�lhe��m.r�T%����K�ez���c�������Z�V���+���aXo�ӑ���[rZ'!E<���8UT�\��̘Y��5tz�?㱞?X^乴d��W��=Ρ~C�j	����g~�/���3L��t�tD�ݸ�Yӌ���H?��қ &�x���H�S߰�e  6َ����$M��n��.2�eX�q���!�$m�f�B�$�,=[�rg~�E ���Nv����f����m$osT�_����w�k["��}+���oS���+ �� �d�QD�ڨ-'c�L��x
�����ۣ�\� Fc�⾛W��UI��P���������Sj0Mqx!������:����Cy�>�/l!+DvU
���`� �t{Xb����̃d�j��};�) 7��/1~���"��`��
�巺Y�aM��|��/;�X0 H�eTBOJj�C�nE�m����>Ps����Q+~Ah�:�Bj	�0k��w���#�*V

��?C�u����m��Wۨ���;?�i?;
3�8ǣ�b������4S�=���t*7����l<�o���q�
�����H�Fq�� ��`/�/S�u#A%��y���)57���4K��m��r������?�EN��Y���+����t���f^X�t�lS�"-�JA��R,�!��A݆Xӿ���gZ|���Sb1E�|�p�J�i+>�F�.#\lFfW� �;:����Yd�o���
W��yJ#�^(��l�6��	�ɷx](�ט9ro�o����	��[<�#q�o���SV2;P�sǿ5�b��AKq�X��C��h(��6�L~�!%�x'������Qʝ
f5W��~��9}�5����l�u�^ĨF`tr^`f�H���W#X {�6�CsM�߂G��V�@���{8yR��@Yx�5�eF�ç�`�LK�o������}��aW2���w��{0#�~KyxZN��J�L^$ݨ!f��f*�٬�(��IhR�����eA|�Ka����2(/AU0':�,���Q0�����[����!n��mr@�x�� U��>l<��i��԰|�Z��@~y�A��]����]1*j�9/��ܼ^t� *K��m]�H��0�θ���T�зj=`t������4��Mz��1&��!U[kk<��fC�W!�>���BI7���Ãtvi�,��(�T]Ɉ�8��g��k�|L���@�����G�Mijk`� ���Y�[m��	W���H��&�>��}���1�@�Q��fy|�h��������V	1���z.�ޭ����x[��n=���<�3is7Rj�^#+[X꿬���4L22��wT;\��Z�օ��q��v�{i�s��QU'��Sן���(s��A�&j�v�s4Q+�S�E����.Ϻ�����@��<�T6�Ī
dy�<�?M?P�h�υ+��Y���C���=}F�d�����I�^>�t
X���q79[2�Y�e1�$F9��Z$��H����r�wi)[>6�z,�b��/�NT����oFV<�b>��8�?◥I�4�Z�����8�}���P[/U�J(�,P�ߍ��|+����rs��Dqx�f�d�T��zZ�9�W�y�y��F�l�
J�.Dì�M7*��( ���$(��`�����W3vwwd2`w��B-���#3q�A�[�?~��6[r�]  �e�T�KK� C;�0�j������������@�Ej�p�f ԌU=����?�p���0�ة'U���[k��̗=Љ<7B��K�W �B|4��8�d�C�[Gh8~��a�\�GC<���9���c�V��o��c���q�)9���M�(Zq� n��9����"SQ��WN�+�T�d�����0X�W�W����Bp k��flc6Ŋ� �v�]��ũ�V�Ns��X�?�x�TrS[�kF��^���LU��..�ȃ
;��=GEKY�����˟��_\}��
3�k�C.�	��Yl5����)�����<2�\q��nx����&�ގaJ�X'u�`�W��c�j�Y$ ��hֱ�Ț���/�X��q޿���J�{vR�`��e���"��bk���.k�F~�McE�3�����V��E�� nt�)�kl�_��ש����Am%9���pdx���sS�����	�yTHE�ߔ�F<6_�5L����U�:S��t1�pɚ8d���)������}��Ctu�b�p=Իb7-���v?���V�_q�F�	���A���
E������g��BD������	���]�M3̚�9~�uo�]���U��Ab$<��M�ޮ~��̭�PpKF���
��?�I+����¬&�ۧ���ޙ���0ֵ5��.X��:�hƃ� �2Z��DA.%�8�M9�"�(q!�|4�⋅t,��[���!�����>A�2���x>=k���A����j���dHF����[�A���G�Q@��ε�}̚5��h�ۥ�����h:��K�.�����W/���R���Õ��[4�9�k�z�Г{c�q]���Q�h�GÙ;�4����� ��-N�?>�����>2r�P���j�7�cT�3�����!�`��M~{J�����i����������<eTPH����;�oh2�,к�@��hZ�FX��b�kݐ9�Y�d�;7��m8��D�Ie=�|E��+��Pz���/!�:W\�ˮ2_��ƻ2�d�����Uͥ�-Y�������Vf��N�kD��;y�ߚt�q����)���]�XKT�*�\)(��X�97�>�>��Cs�5���Swהc��n0X��
�=��	Y��l�k���,�g�Q͞5���T͡4��>��j�c�(׳��>_S2'� �;jg��e>ĺ�]V1��o�֏S?w>k����!�`ꪗEU%�SA�!�ڟ3���o��bq�%����r���KĿ		ct*/Y`h*bD�K�e��=��sQ����c�&o�+�?�$�bc!��Z����g��2�D�d?^�>ar�$�=O"�k!��q�y�G�eL�k�ԡ�X��O}<�\�[�}+L]��=�ک�ۗB-�&�x|���/��p��*.E-�&x���%�hR#����7�k�Z�3���I�jk����k���a���N�$/��8��<,�z*ޚ-�;�>z������$�DN�.����]�F�]V�>	�z�uM4���d:e����%d�������ʝ����� ��-dU�<-&��\�[ ���)�>5%��we���%�r��r��6R���X"Q��@&G�h��x���e\'Y������f�^��BX�8��}n���AjU	�+��r�,1~N����j~Vg��kq>e#�i�����Zc���L�~���O��ޚS� "������"��C�PP �0�=Lm�������uy���\aK�d����Z1`fud�/Q�]�%�;y�#+7�Ҟ�P��n@�$2.r�z��\n��]+��瞅&~'��{pg�a`��RrVs7�]{]=@
X�?!%�>Y&{����;�"8 ��W��rP\ь��z��F�"�eK����`l$� �۟}!������1Nc����E„�U`a�������K!�i=�:�*q	)�S���	� ^r���U������~���HX�f���i����!VI��� �v��7�����&�>�Cu�����7��%Y�s9E���g����nD�h�i�gG�Mj��>�������8F0#ׄ��M��rd]R
y ������}-sA&cla�#<	k=��L��HF�Ƿ���/29l��~���_��g�F�&���6V�rw�B�! Z�� _�"�\:m�W�9a.�����C-4�9��'v�ԃhiKو�����-1�