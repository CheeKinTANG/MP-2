XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Eo؃ڶ�8q�MNZL3#/|[=q�X� �n�s�V�R\����j�g/�<��[P���o�}(_� b�:��W����v>cJ�����&�~͚�qa�o�֓���o��7o�b
_���;eH�lN���K�8�Q��&���0�l3ҷUM�����3|k�{BU��?�T=���OڀFG@gF5�n������+��cGb��ц�Of��hV��6Y�a,RO��`�2r�o�u����P�n�2��]p
2.#8b�zu��_cڰ�e@��.4��e��IEՠ��&K[S��L��\.�|l�{ĲZ���Ѱt����V�8Fs����� �0�=�����n�!�|[�}�l�RşWDCS#����5&ov��Ld>b��xLz��}��+z���G����{�Y[p�<h#@u7����ݐ�X�w��"Yl5�{��7�W��}�Q�|�[S�f!�W�_p��[�8��\:�6FZIF�����{��W�K���!j2��P �u�Ú�ai���N^��WE\��W :f��$��������p]���&|^Y�^�t��Y��A`r�凲�ɝ��/�Hl�W�ِ��3p����zn&]16�8���cE&�ʶ襉9b����&��(�x���dH��X�ؿ]��ǜ���]�@o`��:��+e�&�����y�[8ǌc���0��n@(-�q�0?� ]W�ӯs{��G��?/n�B��}��UKsV��Q�X{����T�����XlxVHYEB    3e93    10b0k�Fl���x��-�w:ЖVA�C�߹�3�5ek1��[�?����� �k$��ï#�٠ۛ��=���N�����&�x�l6�Q���qx���-7�w^�TW�S���,��i����ףj�Hڲ���	�C5	d%��L �D�M:�A45r#��5ˠS@ܧ|՛�W�Y�z���]�+��E$re������`6�wả3ux{����TѦ�t��;����Յ�a`Bg��AH-�L����y܄=���J����Ww\A5W�N�b9>��Q����f��qV�̰�\؂{�.�Q�%�� p8G̶�1ћY�/od��R�����s:7���w��=7p���٢f��"R������H��~}˥��ٽ�����Ha�U��4�� ,~W,�m�R�����$�D��\���.�}ug�y�&��g;�������3�&�<������L�k������O�5�J�Հ�Hsh|�o���
�H;3�*��K�t��79?����|l~��;�%��Ý�?�Z]�|�Cߜmn�љTF"��cҋ��2L&`���?��$�z��?_#��]0�(�gB����޿�������i3�AFZ�J���|��lm�)u�Z�n3����>��sB��*��7���?�)��Pd���<�.1�Ԃ���7e�ȟ.�w�����A����!wE��Dd�w�5|��������O#�1r�#n糮?��w���͂�q� ՊöQ�Y�7w7�t��Hd���G����]3�Y�P';0MX 5�S�t���jl����eiN<j��a���a�1c�p-��Gd��Կ@qh%.m�:��N������L$�Wt���[��,hH+=����@� t�B�|�|VPO�zbB<��ۈ�\^$n����zȘ���aL�8��DLՑV,<��خW�#fK_�e)��d��-��:�O�{
��m���M�T��?�+��O�ԕ���%�� 6DY����b���>��0,���`�TI����)<f>�����t�ع_-Y�俻����H+qH�+uc-����n�lE�k�i,�i�D5%Z�t�7Oe�?E--C�;fW�M<{�ԏiѵ�	k7b��\��ӠtLO�s��_�h�sX��Jâ�v�b<e�����xZҀ��
����A�STx�f���)&z�ٓO��4�l��=�v |Ѹ�r�~3}L�ZOm-r�2�����?�W/���)�Rܵ�-`43�l���%	��F���+$B,p�����v�򓩔
� �A����d�ƛ��$�:՜z(R�.�,i��9�`u�v ��U*�� \G��}[�F����VM%1��8�M�'V�yvq���R���5P�Z��g�ڍV��Q�{� ң����3��duH�m�4G4�x쫉�\$x#�b*�!m2mZ���Z���3������D�Ryt��O�t�k�}ܪ$!�t��� bq:�HE�g��5��Y%}��/��Fw^�j�~@���yqL�چ���sDi��y�!ٮ�ೂ��6�yTf4�1���)��[�c��x���+���U5Z�J��EL.^��S�|x��o>��Û[o�i3LQ�`��=.|I��v��Aٷ�7�e�$�G��p]��.Z<�����D����<��=qP���Q�/}6������yI���p΄�\�"|�C�^7P��y`|�PnHQ[���|\�e���-#�	���Q��. @k
' w���#����U9�4PP��~<^)�h������=E���!Y�)L�g>�u��R&I�lȫ�<����@����dUN� j�	����e���{_�uMݳ��[�H�vn�J3�����r�Q[)>9�w;��U����7�$�-�d;ޑ����h+<TsXZ]�#%�J��-��X��'	٪t�<��5�V��M3b�-�+�0�dt&��p���+ԑYT������Z�PY̅��p�a�	�e�m�~��v��UM�f��jG�n�~%�lٗ�':���D �Z)mO������7�N_Q<���.��u~�o�����ul�	��M}G��_ܽF�q�� jj+�J)���](Ŗ����^��U8��JN^�����7��	��[J(Z �/Ϣ�;�xY����z*��pDK� ;���2�s)ϙ�����.�aq ��\�<hkDPQ�#@A靖�����qu1�xu5r��[�W��>ʴ����I��G'� O�@
Nv����� [:�
���J c埽�Bʹ;EL���S���Y9�������Lԩ��<��,����ߌ
�{�-���=sT�P+� Е��\,b�Oj�$b�F��k{�u���W��1:U�%?��[2�=yؚ�!�ceU�Fg�>W�#F���7\�&%�q��̬�5l� �I�S�dj8p��A����:��~�Ӗ�U��*��X���o�%�C3�͚��\sKMQ&2h8ޫ��3�~���\��&9�p*���3RJ!��<�jjС��,�(`�g}��MLGG�YO1��m*�ݤx�$���S -4z?�͒[wr�Nrd3��'3�-&9ǌT��Ƚ�I�K8��׻��0g��#tk�צ�L���ǳ�q�5�t�~���H��V��U��_�O�Y������S��WمV���JUy{xL�L3>کuU���b[��4[���Q���#+[�l�ִ7����Ѿ@�����{����?�Ѩ��̧7TE��0�� @��T�"Q���_I�菩��}S4gV�k6Gn�z�#5zO��P��@�~j6�v���޺�ʚG�Zj�N��/�b���;V����Ѽڙ	�*���<l~�=ŋפ70Z�"a��X|�h�2��%N�@��*B�|�T���>H��#�B��e��-&�S����{u��Ma?��VP�v��2z�UIw�}����qH��dζ��ܼk�����D�_�$O��^/���D:#�0�|�F�\ ��mD�?��xD�684��0`���p��M��w�`��(b&�>U_�y.-Baj�e�����T����GO�˰��CzF�$Ş�F���{ަ�]�	���[u���K�:x�\Fk�&~�9虶�q�"3,�M�0G�o���x���ңǖ�;
�J�$(�l� X�iIT����O�0ƕ�K�����HV7�����"�ݣ��Jq'�j�����@�"
�>���j��$Ϗru��NW����83R����-y���NV"Aq߱�av���ӽWG��������Y+
p����������k�q��s�a	ޚ}�-q�h�F\[�ë�d�fr��?³/3���$6R�b�z��Hsö5���3�A[�@[�2OJ��g���b��nXy��b�'ɵӭeO Oz��228$�!#(y�8�K��'؟�M}���E�"X�Dn���b������C�4�bX����9�]�7iC�`B�&����9��x��Z��#�n;��%T6!�3u:�����T���j��j�ƱA�4A٬�&f�}m�����eo��˱���t���6�u�E�Ƈfm�o��Q���� +[�/��4Xd�ˢ����V��C)db������J<EL��};+�Ԫ=�����f~��'�/���k��S���F��e�G�n�'�;�=�S�o !*��/MG�Zc���!}4=hB�P9���#BP����ɌJ��.Fݼ\���"��?�Kr��G3�g��W�``��7.����Rs��"�I!Q���R-k�"���(}���
��6��6�z���m$�Wy�� ����1m<�>ei=��I�D��dV٪p�PP�ø��eL0��맷k��M��v�C�K�#Lj,-������'����n�c�������\?j�	�KI~G��̹ܲK��.��R���Fz���d���$�>��y�����4���}M^W��S������#6ix�SA�2��o�������d����%ݨ>�����l*�C�T������Q}���e���b�P�!n�4��_�nxڴ]b�[+X$�$ �(�$��?�#�%K�Pxe�Ew�����9:�����a׾����ǈ:J(��;'���Gog����*��F�j���{dL�~r�-	:%s_����|T��1x�Z���^�7bRg갴��>��靖�"�s�<���9 R��`�x�4�'�~�6�U/|�EJ����'�W�*I�I���(