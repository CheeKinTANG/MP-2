XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g,�}�����;1�1�)�خ~�o�)!��eL{��|�e�әG(H�M}�$��]�/9�h�z1�Q���r�����Xo�zihN/2�0�D�!�k�s l/� ���K�
�l*��V�}��ylm��-�<��wW섴�������8l��|�=[H�Fd!~Иx�z����v�{��!Y�>���ۿ�QFsLe�G�x�n�{��x �EK��b��J�qH�N���KFi��S�O�֕��Ϳ퉨(�WJ �Q�M��1H���}�{!��6�uW5,����cZ��nNfG��?�a����y)�`��g�����r���)�4�E��WX���3���򅍤��j��]&GI<2�Ъ9�%OG�H��Г�,�e��x��l�t+��ѡ���&M�ҘEx��*~M�)fb�}i8ƿ�-\�4>"8BJRБ�סS�W���M@��N��+�M�0��p�(>Xx��tV18����3�#��	�x�@���%����Ε[�r@;Bn����T��6uc��0"gّB�H��`��H.��t��_�>f1�|�{[x��\���\�==�Ǿ��Q�;�
��Lm6������DVg�A�nj	��P4	0���s�$��(N#g�s'O�Dq��G��p�~�ϒ)cd���f�e͓~}�i�&|g"�8ׄ���t=�uA��_h�{���X�Bѧ�u���t"݄��#蜼y������ĥ'�o�P�%T�nb�0Լ!��/U�y� mzh��lpƮXlxVHYEB    b087    2540q.��lA�g�u���0��c�� ���o ^ř�7�O��5f>���ǝ0%���ja�:=7+��Aw�a��#I�u��s��[���M�d����dd�"��WF�j�ZO�46a>pyd�ι����Q鲣��b����8�+6��G��0�N�E���[,��ǥT��Q^�ٟI�����b
��6���d��o۰n��Ld ��d1
+!/ʕOfH���g����U��w�B���9��I1}KhD��u�F��Ɨ��]�c$�VV��A��üXh�JR�稉h�����U�ա!���Ul�������?[-7�)����.�<v����=
�_���:�vkLm�kT0��5���Ue�x�|�	�\l���X��}��]�9y�Bz/ы��|e����E�$���<���4[�Q�UD��[1����C�d�a[�05�0��f��S��7�)!1�����DO�h�nK�=g�٬7:��������.�<qVe���MT�������~;�,,
`��tU0���� �iyH8lJt5=�zk�\��LN��#z�E?�nͰr7b8G�k��o�X��]X�3l#��x�5��m+���֢�X�7 U�x���ִ͚'f%}r���완��ۆ�%���E��o%ȴ��#��O����'3D�t�;X����>�p�+�X��ˢ�Ρ+����o֤b��y��W�kX2-��;���HyO���٫���&� ;q�)�.l���^A~~��4��j���"�zD�+a|��l�4Eظ��&!�&�
*����A�X*C�8�l�hÌ<�V�,a�L����#tN��ގ�q���\�@�?m� |��0 ^�匉��5k�6ڈ��4�~�B"���� 𺦗��� U|L�*��D�;Ǘ~֛R�F�OO�q]�ɼ�/ln�t��$ޫC���`�m뇊�?ao�ꪏ�f�A�IȂ��/���zTd�vY������3sy�wM�4����8�+t�ƵLQ�>r���g��n�w��*O8��O�U��U�\�& �݆�­p�;,��a�d��_P_H�"�Ʊ��k?m� ,��bLz�[���e5L�y��|�x-�b������兪��~���� K�8�J��kF����x��@�O��Dj3����J�C�&Kv^3�;�(���5�^u��o�k��-�������4��<+�$�T��߆��F��9�d�P����8.��~������8 �
8�
)m<�[,gv�M��$c	Ng7�(�L�N�WJ���Qy�dx����}������q�=�~Q98ߓh=���T�*7F�׭�<���.�? K�.G�K�(.��a˳S�f${a#jƖ$��u���{�����T�)������Լ%g�T�^F5T�^4�{�l9G�ǌ\V�]5��wi�6b0@����m��c$@怣�q�fRq��c��/A2�IH3l;�z�C�� �z�Ԑ����a����j`P=Ϩ��Jd������4n�f��6w�ɐ"��ٵ����K]�B�o�>�pm���UZ� �:�xBB
@�g��(Qv�8��.w) ����f�D�kD�1�qR����lNj��i�~�қLq�0'
~d��b�^�X����jlC�B��Į�߭�պ)�g���ґ��b�j=����LQch=zg��Ԫ�wd�+%�܀�B�`�����4�
���+b��cJ���.Ш#y�Z��h�E!���ln���>�\F9к�[h� &~�&�B����R"%���R��������>ڪ�`�T/\^�uey�eL�a��P$W��X�@6��FL� 4����?�#Q�9�`��]�(tBY��<��U�M�A�9H.?��ޤ#����E�x4�`�� 0�"|V�$�$0'�lu�U��;ޱN��.m�|��S��QUR�e����,.F�}-�� ɨS��4�n���֚ �����`��Ts�,�����φlSc��jn��KS}_³�\> ��7@�7-Of�
�?��p#��E���ɐ���@?။�MՉ�v�9&V#dD��ǆy���@�[��^E�
���5*���-�;�J�?�y��.��K=P�O��Ụs'��= �]���H�j��*>�7U䬴}d5#{�A�<����)��WP�I����jYp�Z㽸���U)eu�D��$*Mn'��}�JE�@%-�E�A�=DH��?6�4vۉ��:=_C��u{�\�pEG�zq���)��/��v����U�,��g	��ĩ3y�n�!��A��x��;pԉ������.�2���o�#ԩK�0K�t2 dQK����ƛ�tv]�b��+�XU2�i��j�	3��T)uc|��-k�x��w�d^��B0�l�D{p蠞��j�+�*
,)'I�?jlR�1��e�6�'7�)z�����y`ဵ=���TP�(��~w��D
��R.'w�Nl"
��M^,�;ѧ�c���V\����4����uS�uZ�͑=���`kD�>�C��߽��@����c�7C�h��3��4MC���V�l�������nJ?���)��K<�,���%{������������+�1�i��݀��ݰ��d���|V��x��2���}2�k���̟O��L��R5��ʷCS�hV"%��,L��-�����ZGn���Y `bS�J�6EC��!�B�t�ͷ�h{��'�=�'��*C�l�'�U>-��tu��J����&	n8ZkH�=7�;Z��o1pQC~���6���\�W1GW��t�N�zލ$��	�~I'�_y ׬���%���MlC(�-ƣ2'���/%�Qt��'._Jdx�"�!�+;&��V�8���`�@6�A��f��_�5�����ۡiy��y�Fh](��5$}q���.f"ǒ���!�2in�+�<y�@�e�OR$(\vU���o~�㑥�1�S׆����I�g���Hu�a
rkd�7��W���O�Jn(.􀠯EN���2W����l�G��x�߿��1f��Χ����;�O�e��Q�O5�Z���[_A�p�V��C� ���6-Bvw�����`���U�Z��x�*?9Sx���v��Y���$: �'�Rp�#h��$�!m��a׺ƪ��_Y�+�+�C���<�LZ�]����� ��W��?��^��{�H(C�<@��<���A~/X_<yS�[�.:�@�1���VE5������D}�Dp��
�YwZ�Ar�ө9���>����RƲ;jg�ˢɟ�^@tz|��hn�+㢡����v�Y�W��&)cG=�%#wJ,sT�v��/�5�*:J��(�n�z�n�����z\�V�.����NJ厺������v5��a)s�X�HT5`f�V?�����,pLYF��_1X�z���!�;�2���Y��]�)lOp�b�7V�s@cS��XD���
q��V��rW������;�l�R2"6;�-����6�R{q;��>�2L�@���NxzL"�sCIy�c��qv�	�q��Z���{Ba�c=�h- �gn�K9?tm��7���Mkqg���Biy��@�(������D�d\U'���0{K���0�q�$Q������e�I'�k��2�3�e��-�݆JV����S�%G���^�=����ͪ�z�(*��4�Z�%:�����9P��t���HP-��:�K���dČ�[*AC�Z����#P�1�s:�v�.?�����\���z�)��+�i�`�������^�\)	�n��#�V*��9̩�z���;�!�{vG5 ��tf؛øeǒ���Y�{,?tGwb�oc5��V�	���=G�{S{�|I�\�;�g�ڨ���K�<��#��c'�q.Rn@�f�1��+�7�X�4�0����_�=�;Q��Q�ix`�HU�]T�j��7A�+:���V���.}�r
�o��2S ��|.X��i���6�\�r�<	қ��e?e+�:_����)��������;t�o`�=�����$w���$��IN˄�Sw�;�Оb|�	�6cJ؅/�ȫ�X6q�rz>Q!�N���sG�>�x�&F&;�����X���~f;�a��\,D\���`<�j?8�Q��^ʎK�
VL�k؛�D�l��b����4�Ⱦ�w�q�Y6Yɰ�Hi��������d��3���|H_���5�	T�\���I+~�� K�5��^Ѐ��UQ��y�WiD43�Tt�5���@��-��
�+��{z�_����
]X��^�[°,D���0�� (Z#��[�ۨ�,H�&��C����T�2�"�����JUn3MBB;+RT6!M����Z�h��a*�����u),�1P;ݛ��M,���=[Z��w�z ~�GfoN!ģh��%�5�M��)|~4&xCZ�>��7J��*���p�����cQ$%�`JVw%SQ�G���u���u���
�9����1}d]��k��7�O�x���ɉ+��T��L9�P�ȗ��Bwq}��:X��`�Ւ����X.�c%)J�;O�g�0�״g5����&��i#u%/�{|;�T�T��	�	d�^�'�h��[E��A؁A������ɜ���V�y���(I��z�E�_�$ ���.C䔤XY�fN�8)zUN���5<��Ӽ,b�I��Pkf�� 餍�BT���0α��n01��)'eRn��H���(�"@Rf.a
|��b*8}?ՓW�G����I�k@p�%=����� ��G,����c�9N*޹굍��z���jS���$6��������:�6Wd�,z)BM�3qS���z�;��]�O���O�d�wB�:��ud�7�Nɋ?�qZ�F�����B6$�K���ڒ��#���S~Y��ן#,Cu�y����<,=u �-��k�x���<�]���_kQ��a�f��=;B*#1���+:�[[/���jH���[å(^���43.]��*�[���	�V�11'�ծ9��L�vR>?=��(��X�.��Lx�i����WY���Pe�.J,��@��I�I���޵���2�Gncff�����X�$�t�r�X]��Ɠ;�1+lF��r�~�q1$I�WpD{�&���iG=%+���%����G<����N�/�>o��Fhp`���f>�ưU� ��M�䤕H��)EԱt�^��`�N�R��Y�7�|,,�f��na����Onw��H]��*_Z�4�1�/�0*o|�ǇЇӃx�=�R�$�$���VD�����Ȉk�KEm�Y{R��Ŵ�������Lʃ�e½eF�u=9��{1&Y��8Kɞ�2���|'���E�#����?�X��"R�����ـy�2��$Y�Ƒôۻ"ԟ���ߖ�Qk>�@���?��h�қf_��V3��$+�.��u�w���LY"��Ҽq��g��^lNc��4֖e�n�.�Z.��\��f�J��Ż��
����E�b�?	�t\��H{Y�K�S+�����%4r��Y��1���'�Z���.��� [�ۨõ$����A�s�k�*趵ΈYޞ����E�U���~qe�y7c2���(��v�e�zj�E�%f.h�7,��`���}�(��]�f��c^��	���R��>/M�pJl��g胖���.��J	!{^7	J�OZ���U�"��,Q�I��
zrB���N�\D�	��1A��t�K��5NH��+[xq�e�S\'�����e��P��=�� ��U�M�@}Rm2|a��$ϔ͗���9C=�Ȣ[U}ե�����WH�'��>�����&��5��
L�ZFj�}dW�ޘ�e�Km���R%������"���Ʃ���UfyB��'Õ�m��$���V->eN�����n����6룤�@�n����)� Y�mZT� &J$��\�`跧�N�e2�"4��5�xL,���?����5�3 m�
����L:�!c��lw�E�fFB��M:�k���(]V�X��Ķ�$Z�0B��~I1�	^ɗ�z�\ٍvN� �o��u��2&�m����k.[����F����ô�S�]��|2
���E�p*½��77z��!?S(����ӎ}01~g�?h5�\�P���d�,���h7ِ2���n�V��R��.�Ve�� �EOq�x����|��=Y�<:���,�l�!f�´x�~��E�5\��A�1N̕f�_{�f������%W%}�)��j����;�Y��{'yUs��b*�`��$�wX�j�h��i �e��	�n�8_M��Ԇ�^z���%*��k���Y�>f��͂�)�Jҳ�;6��2�	)�k\bzQ��}���#�)���-�k�8�B��q��WT&��:kVf�[�gw��=4;,��!s���Vmy��밐����)!�L_�{0��
�����C��HӢ���{�h���Ѩ~/$H
���Q�gZ+���4٥>x<��b��d�����b��O`3e�*�HAJx/��%�o{|��y3#�c��t��j�q9rW��^5�,��	쒘Ri�ta�@�mej3/)J�P�� �ŴYc� ��>�[+X��ra�ֶ�՟�XU掃�гY��,gY����z�c��(>�����60��d�RtTo:vs��YeY���W�"�RZ�ق�4g�3��Jm�Ϣ��h���g���N{�w�k!L^�DϹw	�T h��;
��O��K�*Fd-�c=��lċ�ת���'�|��B��;2��9��_MP%D�8WH�8쯋�X�TNUH�52w��(Ǿ����s^{w�y��M�7��3�az��`#��/�m�xY��CehM���2�����Q=��dZa�1��p�f�r��z��{��_em@z!pw��bK�L�Nv��\ʕ����5��m���E�4�D�E?%�JO�Xe1�_]�U�8�|K�,�d�4�n����gxR����V�g�jU|�A4��L�Ŗ���T=#f��
`��+/M�'�|#��cEDS�距����������E��35� ��7�����|}�<%���u�]n΀	&;�jI�ؾ��*�L��k��ƪ���{h��Q=�di�L����������UA���e2>��S����N5����N�������A�O�d+G�8r�}�;˳��� 7�I��5K����գ�m�q�A�f���d��g��/�u�1�B)���:���T��Ϥrv9͞ q�cʣ�׃N��H��g� q1^�*�@J�w�j��x��H�*�.��w!�����i2&�G{m�� }9&F��t�=�� R'�� w􌮎�4c��Ȼ��1��i;Ȳ�{$pF�����կ�Dt�ZG�qP$[��W.����܌\t�&'����LH�H@Y�8�L��N�����B1�TS�vHh-�9�'�enVT�c�#��bQ�C�P�t���v�|�� �v�ZfPZ�x��=C�I�t7�)�/os�β8�NOMV��96���q>ŝ�Ƙhq��d|8ۜ�s[k�l<-�5z�{*�]������y�"×�� ;�6��`T�t�8�dm]��#�p˺�&�jעi]'��8�_���[>�+��߲mx��)������۠6UJ@!������!Ji�E���!���é�����%M��L ����� ���>��_G4��Z?�W��[ȑ���zF@�Z�ܰ �Z=ȁ���"�����54Id�5��P@�~�<���){�[E_dC�ǽ��LRnR{��0���7qÀ��`Y�iP�.]p�S5���P�~(as]��? ���6Ι��\�|���V}��=R�����3�J^��ې�6Ml�a��ċ/B=���B~zc���1��E�,���(]��� W:U\������XՍ�j֚V��V
��q})�$^���-u��[�i�]ė��I��2�0H`wQ5�GQ|�
��Ue��j��n����!n��i������w
������
w��TLˌfA;n��q1�Rs|B�l���س}�N�:�v��X�@$��#��X����1!K���z߰9I1.������k�`�Ϊ?�D���ow�$���B��W�m9*'��ל��"�ʐ�s��ȍ���FՊ(b�d]�zg��Gۋ�]n�R���2hC݂��S���^��dR�m�����!=8�a>;��I��Pl͙b+�0���3Yq��BR��u�&f�]�����֊�bzY�g�hT։ZP&�2��65h�	�;�Vq��1�|�Y��9�0���س����UV�$	����׀K���9В����^Cd��'��U��4���ٮ��&.p=�ݶPG@n�%9XlT�n�#����pS�}tf~:*Zۇ	n�`p�rf�?����n|k�B+�H:_G(B.��_ eq�����\�,d�?E����٬�郬�(�6����ŮW��e�}},�=��CB�Q��V���cr��~�6���~�/︂q�3g�O�u�m�ښ�a���̗�� ����ZU��M�[f���n��Z��C����3l��d�)�R���~�Gެ�w�NGG���̇戥�x?�u=��(]��@���q�2�U�����-�w]<�'~���Y�e�RB��q�/(u�Vd"��  ��Y��g�v�:S��ER����G��6��c��(V��K�}�,�`E�/"zB��:ȣ�8�SSRv��3DM!���(���<��}e nO���B�|��=����b���]��/Z�N��8����_	@������c�y���S�}%��6Nz��Ǳc�7�#��i^���x�s�);y���TN��߹���.o��V����t�)u��]5}3R���`��v������v�C�'hO��.\yp�$@��|���B�7k _yŲG�n�^oc���Y�F��2�U*��{���2HA99+�.��v�+L����G"�R;�e�;L%\�ޥT#��n7˳�/}��Sq�+�ڗ�C��r�l�Bp�I�S+�U����`������?s�y}�N3��I�����z{`��R�ໃg�]| ͵	I���F�ˣ�2zY�oq�_ĠE�$��-�n/���0�$�S�|�"����(��|���w ~ ��:�g"��{��;�j�Mi���8L+*��E�78N�Q� s�L�3n+�9���En�h4T~t:�N��M��煡+��g��CX��な��A3����T�՚�_��2 �I�-���ԍEկR��:ހ�8�u�n���I5�J&���{�h�	�a�(�|�s���i��lݕkk�-6w@���G��߱{2#BU�kG�?�]�U�vD��z�ƪ��ئA6�ߙ#�MX+]���