XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����rh���L^�z�'�U��y)��z-������N3���O���Q��sM��$�d
�×H�-c��·y��}H�_$M;��>"A��.�U�&fw	��pPїd�Ϩɐ�Z������Q�Z��ն��CŸ��Ԝ7�� `���W�~j�vjU񊄄�����<
�L���'oֳ��Է�UX7�@�kȴ_�/�k�SC>L?������U���S��Ǜ�%f�G��3 H���}x��bղ�z�W[���S�ڥy�~֓1j�ܗ��հ�YX惋���褧�}ĸ[����[�sJ@F�a�T�
#�����ˀ!�_сO�*m۾��I�}����l���J�� j����+� ��4�
�m���%�7�D�� �m�O<��S:�2R�c������x?����V+�z#U����4�ҋ������7x�c�&JE�5�bQ��^�dG(����|�*�tY{m�5Q����G�9mbE̙J��~�8���ٹ�p?݄Jb����9�H�4e^��&4s� ��ĵk|�	 tb�J��q,M@�ʶzd�m��!����+��u��H���?�$Rl��~��0#�.�k��5Ɓ��C��Jn�^SY2��z�zU>����Ȉ���3z�H炢�����pƕx��=Z��ry�J�!�f�B^a)NzڸGd��M����x繙K����6ģ#"*�7����փ�u?�����Wo���eƿ|���&o�$�<ˏ�Ue���˓�{3���XlxVHYEB     e07     680�d�|�o�XN�OL	�1օ�L�)�5a$&����sM<�?��c"e2�����BHK��8�%�#���$�c-����0�6إ�wQhx������j�p����S��k���0.*l�a�����P a���^X^�� ӞLQ��"?�M�Щ���Ad,�\}2O���@;G �c�=��T*Ӏ��p8�d�j��肈����������ʁC¢+o2�P*}�B�@����М<:2+�^'�V�
@�����0������sD�Ԧ��+��ad&�C�� 4�b�q^$��k�*m�2~�N���w�$x��O�[e��w1)����,�)m>t:&)l��9���Pw}�������XfÞ�b������y畝�?�,�����"SYQ����zǥL�YS������ѝ2§'�Tڥ�S�W%����÷Sޘ�PT�/��w�Z�Hl)�����$�]��z[�y�]�_�T9Z�$v�/C�|m����ym
0��j+r��31�	�t��^;�7��(�^��O�����S���|�4�=�6�^�Q�	�|:�!!z�S;@�TL�w�vYe(@��e��)�E3$�N�*���c��ɜ��'��0y�Y`��*C����z$>�>��2zhV�;[$:О�/�*���A���9NM��p���_{%:T��._��,ĀU󾶉eO*���"'{U��<�["Z�+��st$~s��p*��d�2%�A�z	d<�:	٤L����H�s߮Xhf p[����x�0�9i5p���\Z�3��7@������&�抠
�Pbu^w�jp������jӢ'8��_�'�I��4�$�J9���4��/t�� 1���C[�9��%��J5��[��y�Ė���!��}��¡=��PDg�>)Ce^N���!��h�#r�y�����W�=�LEVqpJ�	�p���ΧB:� ��b��c�H�85ɹ���G�ZH���,P�H�0���c��Jv���!�gs6���B�AU�@A��*ir�G.���`���������mY��a���7R�s�]�W�K!��K7�bϜ���ݛB _|��#��X
�n�E��z��~7�,*�vVﶯ��C6��9���h�W�BY�O��1��A_'� ������)�r��,��bd���+w+=��ݯՈv�K���z=���42-�EڏD���sGI�\�x��[��"?��c����f3��������k{�#� �q���<�j�P���*��-����|�x�~_I�4!�FS�A���ù��h��j|_��D
B�SU�g�C?Lտ���7�9�/Üx����C�@PC�4?]����M��
g
z�����-兝�:��|v
�U�T2�g3��"/#f���S%��%k���٦�]@��bX�d����!d/Z����pB�~��/.�z/h��	��T���^B�z�?�{�#�D��K�\�B�3��%a^��m�*�-Bg��e�-S�����OD�*� e��i#�^����v�C�ۻ��"�r�\�w�z_��| �9���*陳F�{��n+Sܤd$����5}"�*pD��Hf����Yɋ\����M?rr_Բ)��1���n �G>p��,l�ʟ����