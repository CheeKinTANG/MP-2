XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F��(;!3��u�g#����[,תn�DJ?�,7��p8��	�z5k�ǋ�'�����T��þ�Hh�@n�N���KOYO��I�v¿�Pyu�^&�3e]e������<|�R�5�[�\�jo�#c�i�@,�@��-��~�� �kٸ�,-��7����U�����$e�)�N��Qה���.�Ǥw'�Z�o&W���T�S�ۭ~�C���ͯo"���n��(��P�q��F��(z_I�vg|^��^,�nBr4���gm^�[���ړ{�2T������OQZ%���6�<5�0�>2��q%���h�����0�o�Za��P��<�P�1�T�Aoe�wO#Lf���a���'�pQ��n{�"���sZ+ʃD��|��w��rPrd_�bm��9�@�)�������Cf�(S���s�|Վ�>�������[��������p�=!U(��������]��i�A�)��ٟr_8��"��t��V�&V?�����a
\�ӻ�'�.l�a�ZW0U��~��h����
��*J�A$�E����|[x埄����ŉ����Mk��D��d�]��`R���@���*uz1&L��\]	IL�ıF�(vrW�A�+6J]�	)��/[�6*{�m�e+Q���yR��?Wnб�&S�)�yɐ��yy��@"D�u�n�>HK�0�����,ڵQ}ş��!d�J�\���2�f�3��f"<;~�Pu�%&b0���)��[��f�IM��N�zK�XlxVHYEB    5fea    1830��.���(�2@y�x�(�+���u�t�/�h���7����J�����	�V�v\�<!�
i�*�i�t�&��Ἆg���0�i��8�%s�{��U��~�䮋�	�z�-2̸Qru&i ���F��o��i[����n�M���[sP9�橂�Љn�{r���Y����I�y��1�L�5V�ü���:D��S�`Sg[2�<֯�k��ex������U��Q���Կ�b&;�&P�&D��$�� ��G�c�]q����P�&�w���wx��qLw4�!���l ��aL@�k�vH��c3�vף�J�k�^���%����ߒ���_3�sB�3�DA���8>8�;��0m��
��r��K�	���4��G�X��LK^'��G���>$Iv�F�bCƆ��]�YZ��L�(����B� ��h0����i�BT�������w��1C��X޸��PLkE���(z��|#&�
�L�+��	]ϛ���\��Fl+v��R-0!����y����>�k�>��ن`|��d,�)��º��.���GӢpR�t-i�v/��eH��C_�ZlU�D��
A��0���{��.�%:���5����s�����j;�3�i��N���P�I�f쾿�ߵ������5�k�UY�����:��x�s�����q���*�.4&�W��_���	�R�p	��i�BHʿ��z[�[��L�S �3�&�Dv�r\D�@��9��ҷ�����9Gˍ��������񏠊�Pv�&"����D"��Zv_����#bۢuI�z�9����;{%��+_��ί_�T{�nTd.�R�t'�Ƅ������gw�P���9��pz�s�@x _��_.���M�;1�X�K�V/��=;2Q�a6���eƖ�>T�g܆9j��� F��â��.�vj}����ŖyV>b�0�ن_�X�0>ќN��{��"s��bxs�����Ǡ�/5H0�,�~�;(]��f^���"���V~���că���$��9�� ���*A������3�����4�݋(}ڭ`ZSʮY=^C"���W̱"~�A�Nn���j���t�g0���Ð���N���R|�R��C�Y�Q*���Bt���E=v��(eY����}[/?׀��R�f��0�G���5�^ߍ�M��ҏ�BԌC Tg�h��<R�ioirt#M�v1t+��O�Z���W|i��l+d����V���1���F�c�
'�S1�x�$�&�z�إ��s䷵����xލ-45�����vG��ٵW���è78���}fp�PSX:l9�$ؑ�*��v�o��	�l�9��e��z�7�<$e�g�÷��e�?��Q�ơT��ב:��R�a�,��O�
]ɞ�?(<�u�#W+��V�`%�]�͎>�d�s�����a`�^q����b�'4�*m����}N�
�t�ٹ��� #W��WӾ��-j4�L2�����wb��h����{,��F3;Y}�G�b^����~V���;� �.Oԁ�A����J�ǲ���)꟪��6�x+��zr�R�ʓ�u��f�\�&Ӝ�I��0��b7�<�E
w���e1��K`��k� �"�$�8�(\�4B�\j9����5�tD���l7��5��0×���-�5'lw`$aFn�^���ނ�g+��ַ�����:�4�`�b�1�} dOn*�X�Ud��P���o4D�۱_R^Lܶ@�*�ק��F�v")mCFమ(%�j��p�i�a�����ѥ��*-u���I_�U�}�k��w�E��mG���
>GG�{[?�gl�p��hB^�x�r����K�u��E:>IVl�lE�GۺFq��ӌ��I�m߈z��,����;��;J� ��M}�S�+f畯���!�&������D�C~H����%|�_��I�D&�o9��]/�Ba�/���*�q����С�1���]���_꼒�X�w����?{�����l-îx��M�B�"�_�S&�n��Ψ1��o���d.$��i�Z�W��Z�n���]s)ݥo�Ї�0֚���47D{����B�?�u�.	M)�M�"�DmE��g�:1�M�׹#,x�`#.��M)��G�?��67�C֊R�fs�F�^O��ƹ#�ۆ�*���=�.*2 l�,�YGq¶w�;)��!�q�X/Q{�TH.��L��z��5���{Ǻ�cn����ŅV_�,[`owV������� ��+�h:EX�F͸����1�y�̆/��� HM*m���QI|�0�L'�?�DJ��Һ���x4}��t.בW*�?ۻ��=�*ni���;Gs�k	���D�^�y)���x��UT�b�%hiӞټ�;Dgm6b�F���+��=�����^`J����\�1rw��D�@A%R���-��j�ك��e��B
G��>Q�-C��r]�u���92�%�!���Y��烯C0�*���5$�TXX�R�����˩%��\�vg*��F,3@^ye��dB��j�>�޾�D�ZȲ�u��x�aW&LN5"i]�]���1 ���2�|��I���:���6l<�s�8�4Z�ټ۱64^�1�����vM�eY!@�R���[��~���!�U$ֶ@��,�%[��L�a�%/��H�";�o��y11^h�,��<XQ�˶�b���p���g`��aC��K�����}�H��U8hԵ�����d���4���j3��������~3�M�!��z�T�+���6��Ӑ�t��NP�E�꿷���*�mQ�N��Y���}��GP�\�=��E�|�FVQ�(�>��%�y��������A7ό�G��$T�U$�i ��TBX��5��Ђ/=�^GaN?�6�� ��M~["�dϻ�јKqE��Na���q[ܴl1��:ho#)��/�f�^�xdMB�k÷���Yq�����vY�us�IJn��t�vY�/����$B�M�(g�Y����e}d�t�yn�:�̾`|/�H�����1}c��
��-�m8�ɪ�a0Ւz��D#�J(2�M��)�_B�
�r�����_E�y🎝Vۜ�=_�4R����˾��}2�������J`�5������Ϲ4�]_	�{��t��K�I���!1l�蒍@��W��}��D"H�A�*.S�R���r�I_L�lI��;"�ȭ����%�M��U�����F�2"Y�*�ޯ�糄��{_k1�1û�mKoQ`f�2��qc<(�!WǗ��=m$<��gO5�xy}1�ϕs,f��5# q�v�(�a��O��T~8��=�m��z���q�h'^�˫+Β�RW{�YP0Q�Bh1�A&~�<���2?k�pq��a�����^����&�o��B��W
5�������6�k����N�2�p��	>R����4nm����ҩ4�yރ6,t<�n'4�e�5T��ي�s� p�"�,H�[^z�%��%H��꿭�:Y,�z6���c�B�(m�5�;>�B=^D�fյ[0�PGm��p(��j���`�°T���vI����:�C���v���+	�L7�
Ci���ʒÿz:����4VB.���#m��'��m$pZ�p+�r��#���-#�I�k�b�3� �y]!w|/��kAs���,N���� OnN[h>�@�z���;z����?����{�������c��.��g�4\�/���,��Š\WF�e���b��gqx*'�F��zX����U�Q�� iʇS��S������S��&�q/4$��)PrI[�@��m�������$��Z��X4��(f-�@���"t[�f�=�i7"�u4�܆/+m���%�T�V����r(�i� ����:^0�~�ܢ�{lX+M&4}�y헌�\�Jh���g�<�:72�E A�z��X�K[,-��j!B�n*	�E�>����pP�@u�dk�iT�� p�B��%�;Ô��}�[�0.ɲl�U� A 
��.�_N��!/A�RV� �2W�(�8�����.��[�4�6��7�#g��Q�c8|o�[%��8Of�8%e;i҂}3n�n�9���o��h'�8��B7܊zq^��t��Nf|/^GS�<��hW]U�Υ9���#�g*1%�tt=��r�G�;��OQ¦�T�A���p
���GD�!��.���Q�b�
b�\��Ya��3�����Ȱ�-P�6���6J��J׹�Px��Ւ�T��Tx�:Ƨ#����N��.A@�,��8~L��Z9�V`��P��f	0e���0�"�`Ő����{��Ԫ�EWX	\�{��8�B!ҹV����gY۔�C33�Ӟknu�e�l�!�2��I��8Q8P� rʮe<��K10Iw�?x�r"�]y	k;�e�����j>r17y���"���<�j+��o  �8h�Q h�Ǻ,!"�G�	����2}��x�X�[?FˇY��t|C��%��@��i�u1j.�ķ�#2`��m�{>��R��'���<Oҗ��7�T����W9_8�C��a�C�I�/ra�3�޽o�Ă��
��zX"�[�|�D�>��Q�Ut�˹��V"��`��c�|���;'���[�	 �k�l��poL�K�p��C�Q���G���υȈ�����ds��M׻̴#y?;P��V�<q�-��b"�ERү!��u��D#�b� �<gL�8�ۻ�>p���͓����j��Y'0�o+���W�i���*M�&+9FΈ;v��|Lk�+/�i~�T�%R!�n��~��}��8�P
a���tC�jD?����o�7;u��������Y8�)�����j**d/�?�e1�R�i��Px���q7G�Y��oM�:�m���:?��K)�Pj�4E>3��V��>i҄mC70�KL�Xܽ`fk'r�[i��N���UK�5ض�@��?���˞ى{kk�� �� �Q@�S�q/x�-J�,X�D�� %Kc_V��;��Z���2��G%��Q��\@;zOGIy\+,�q ��a˄fU-_Q㋹�r�L��+DJ9�� ����u��o��x`�/���).�9�@�[{������o^��J�Y��aI���*�����B�
��������([��h<��G�c���T7VKS:�6: -k��*4���:'%���>�V�(�h�r$�q���o/�N���~�av�l����5�OB9���=t��i�8�z���<j���#�0����q��������4��IAp�Im��Vھ�𫁡���2�@�6����k�	��/Qs��x_��t[g��o2��NCx1�<��WW\S���)Q��z��+��6\�4L�X���t�@h�.�б��7�"eS�e޴|�^Px)/��Z��/vIK,I�?�8O��!��l��SLZE|j�㊖jՄ�������Iٕy�`��g>Xz�9D��zh�*j�p�%5�,�vpQ
LCnd��yf�]�8{JO�{g�D2{N�Řg�_�+k�2�����
"Nͨ�X}��<���0r~����:˸��D�A�\��@����(=uQ�%�[.��F1�mI���/T�mKT���[P�y�0hL���?�>YI���Xs@�C2V�,9�))\"�~��~\��TM��uΰX(�x"�@dj����c/�Q��Y#�F����"��+��N���>�3m���M� c]s��
*�F7�2Y�dP�S���/�O�z��f���@������z!?�7ۺRc�
�}��ֱh���p���I��=P�yC)'��z����b�����3�G��_�r)��z�pE�w�tg�Ҥ�Ԗ荹��c�7t{��F/���o�6�X�s`y_��C��/���������s�:0!���4ᾯPZK�{��?��o����CA�)���߁�H�����d��ۃp�K\�f��K��l���_!N�_DB�ڌ1�;��K����>,De;�I8F$�'v�Y~�:y�ak'�Ծ)�'g���o_�viR���� ���8�t�[a�T_s��'�
M.��y��P�z>5��,��呥��l{	���,?�m�)U3��CRW�+�X�s].X��;�p�<