XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%-�Ȅ��-�T`�DH�T����y�%ߒ-i�ǜ��۟��p�P������EI%�bZ�*^�w+��r��t�dǵ�	��ɻ�7��-@�N�(�A��P�gM!8�rʭx�� )��Q��h��*�I2�R�}h��|<��͏o�a{����+�x���?Z��'���,�dxB���ts�Kv�n.���>K�^����� ��aZR�1��i�e�����6����5e�+�RH#W|��9/o����=U.~:���|ͥ��#��MV�ٞhB���������/n!J�Sn��lQ�3->dR�����Cg����Y12�\+�T�|+�G�5�M}|�ʨBJ���=\��&l�x2��qyGVƓ��]G��
��Y[�k����߱_2��P��	3�Ɏq�-݇L��6\�y+|$z�"���"�"����t��|;)�t�����a�'e����o�I�Q�jα�gAވ�6,H�P�7�Ks���V#ҕ��������c�M�P��<�m_�ax)c۴h�k�=��C��;����'V�9�H-��/R�	l$y��~Y�2��"����e��������b�E�3YM�[.��[��/A����V��k|fk����F\7Ғ�^G��]�x*!	�3/"rF)����O��G���f�Y�Ew6��l�c8�a��ĳ?d����O±�{�"1C��^dw_�x����6��r;��ٮU���8��^Af}�;I-,%}Iΐ���E2��;�]n�
�)*X�XlxVHYEB    5224    1740�f1<��R��ay��޾nÙJ>���ZW:���+�y����l�J����+)�da�i����f�V��c���?��%W��vay�RuI�G)��M�D,J9�������O��'���>���n��,�����M{)Vӈ���^�G� OOT,�?r�=G{;y�;K�����)��(v-0f泙o�%�=,�
���:��ң׌�v5��`����e���'��l��\T-�h.4H7����Oݷܔ��	a 2M��"n腘J����C�	&�w�z�Ա��+|�/a�]|�?�ә&�G�K��S%�W�\�;�F!KEj���&J(�!���ŏ�"�륇�D����L���|L�t�9'd�i�h5�/d(ʸ)�j��&'4,�:C��a
G������6��϶X{v��Cb��ّb(�#r��?ھ_��6�]	���3��jfŒ�4�oZC+ތ���*y%��ct6�P�u��(��d�l�|��]�Wr$5W��7j�0�����[o�ޕ5�����0������ˊ��9o\��_�K�	��F�9T�c\L�u㠝ɻ���~���-��x҈\��?���0*�O��������a��8�=|g�?I�k#�Q-��	=��^;�:��:bjx��3Hx�N�6�M�\�ii�A�@!X{�۸��w�R-v�V�R�G�]����A��{��2��Q���j��PՍ �sԙ���L�M�p0{s��8�̋a���J��7F����ﰳE�e�U���٤؞Ń#<l_;�Gz`z���E������r웶�R�w~#u�3z�#T,E�BjK.<0u:Z0��/>:A�gE`���T��TUK�n垼�aw~���d��[�l
A�q�ۖ��pY�NEa��C�V@}��8�t��fD2�U������uY�rR�@��_���)xV�t.*+�4I����}��ט��J:�*�����]�`O�r�L�ln�����-��%U\%ŶT������Ύ�)�Qu�r�zg�kQ�Q�Ro��;_������d.f"�*�xv�������k�&JQSXl�ʱ�
���oo�h�!��ϟ�4[��Ǝ��F�R;v+�0?���
�,e�&�����ί�pQ��׎<Ptn M�D<���jk�4��&9�jXN�㪖��OZ:p����L)aƈ`^D>���P��cv��@�r�<T�	��g��Y�"��e>a�axv�~�Ǜ�F�|ؗv8uim������v��. $үOkB:#��k,D9���Xt�ҡ�x���%z��ֺ4ũ�H^A ��G�CG���p��ϔm&a�sh�Ov��6�p���fpR�]����������V8r�;|�*�q��hD���T�+g�GE��d�1:������`-ò����z���a������^��g�6��{ՄUYhzV���RǔWmV;-m���0Y`��n��)B�=rX����b1Щ�߻��*�=�-�ܴ�	����v ����SJ�	��u����g���Yǥ�^W"</+h�.���i0�dGI9�:��x��w�(�KI���D�-����̶�3�ur�no^�Mg�ro���I����8F��D��$jj�8��)����:4�l���\���Mفm�R��Տ��z¥�dx�W�CS&�[/g� ��9�9�Or�˵���CI���@{W���Hb�����z�,�E)�ѳ��9���J�t�q��n�/�Y��6�@����\�|��F�g��|֥�b�x��A@|��$�c�iF��6�xz$�܋ g�B+�{"�L8_{�ƙ�f$�ft��E���Y+.>�pi2rh�9S�R�|�Sw$�<��\qh��>`eT��?!l
%�+�i,�1���(��v�x��}_����T���uޟ}
��=!赲.������V��禖�S�_
����Rw����_0(mJp7%>C���b�ps->퓂�g�W���k�/�w�N���a(����5r�drnI5��ȩ�u���xk��l;/��h�2��#l���"�h�=���LTy0����7��ıQ嶙?h��┍�D��2�J�0�8�\Z޹ ��`?�o�8�0F)�6�܁J�P]s���̤ 2��Z=xQ�|�.5��
��o5nn�Q�:���=����T��yt6ݡ��&�M�����ߤ��o?ae�п�3,v)'y^Maj�jS��b������=i�>�?B�RW���7v���ئ=>����*A���,\gq��=�`�ZC�vA�ɋr�ëI�^�vYZQo6�D*�������݋��ly��i��}��?*�kX��ƴ�p��c��J�8��U��_�Ғm��|���{�6�I:��t��%5����d�w�mc�5�M+�/�.�a�F3ıg��K�m�X�M�}�*��r�C�� Z3����ݶ�/�*Wo5��_�k���z�z��\;YfݑS�G�u����0&�b1s��O!�M��@_?1�&�{����:6\��F3+#�e+�dfЕ,-/��b.mƁ�qS�rF]-%:��3;kY�V�V�hE��A4}�*X���a���ݞ��#G,����]8x`��\>1��Ct!眈F���G�gs����!Ok_��I��������w22?s
7
�"�+���u�Hj�Ò�l�T�uqM\�0�f!&�Àx(B߀*!�U�<�)�7�0�.]��i+����qnZX���P�i�k��b���_�9Xe���C�E3T[�6��"�oB#�(��&·�5�jތj�>B�[���6ڃ�V�͸�Ιb�α��X��$�8||y|��/��L�XV��S���rP:&A
q�yԿ���3g�06y˻��.��B\q
��{Ľ�r�jF���X2�W�;'�֜�Q���6"	�X�ؾ��&p�˗4���J{�~#�i�[ �c;	���p�rŻܕyD�`3��\���Eף��~�b�z�{׈�9ï�eiC�w��%k�S�	 �1~F��o�]�������d����n㑜xj�G�RL��4^�:��bqJż9Nnt@�xL]b�w��5���?�&b:>;!f���Z�NQ$^�_A�3dL��¯\�,�7*;?��%O�n�k�� �q	[�����G�w>��ubX�Zc��"�8~0磜�=C��b�)�sE��rs����������H}]҄�?PK�%�#V�`+JT�{O�`8�c�FE�3�q�Jwg\{���l��C���'�p���>��E4/ʽ�����ud#��<��*�y���P�X#^�iG�W��j�|P��n���4��h܄Y� Ф��6�B Bz�z�gg[K��e0؍�T�����Lm: ����	�f[W��m/��N
�(qJR~;)�J&;|�ǒ2c��O��@���tC�z�>m��t�6��[n�۰.W�M�vc�˃E�4���I���8`��g��KP����~-��n�����-�/ѬU���أ:�����CD�W!��I�]��`ΣCb�j��TOρ�K��Md?4S��	�X뉩��Y�����q7?Ut��:���c9�*Rřrҹ�/�@	p�f������gPr/oK�#ې����I���B����{t���7�H7e��L�ٯ��R���qL�nO��"fv\���"�L�%g�I��j�14��6�_V�3Ϧ�R��z_��I�-`j���@��Tc��X�,�H�;k�[��&��EnW��D�g� r-v��%FNZ*7���=��۟�g7�ȝ��΃.BŶ��8�6�eJ���J 񞝞����-Y�_}�I*��9ITLĄ����6�,��٧w7[W�2�~�m/J�+��һl�M�n����Ŵ�oҵ��	|�I��a��0����k�u^�w�d��G�޲K �|���i�I��Hf�½�O����8ùq P 4�S/���t���2�if  ���*��4�w@r�����F�&j�&�Te�ϲ3x�h_^�2��2d�x�"��	�Y��IB��wJ���y������<f`k	�^�qN��{��a{�o���Ó�^څ~&'�Q6�+B%ѧ�Lw���Y_;�5�6�U��B�3ѯ��-��ti'Y��8�{�)L�wk���$�	3K���!��Wx&0
�	�Y�:h��R�KF�D��ӽ�>��ǲ���Gc=�3���_�v��JW�f��1qa[��D��y$�/�i�_~��\2�<�/ǲ��\�H P��k`�_zT�կ��ቶ����<TR�B.�3��߬)Z��L������N����br�3�����>8��
��\Vm���i��3�T9��T���"�t���	�c���T�7�'�P��U0�$�����bh*i�2V0X���J��kIZ�F����n�w�8�L�N0�+i0]n'���&=�N@JB}������sω̗�&!�K����B\�TG&��Jq�pA��C ���.0�wf�JS�׳�px�#=�X|���M���?�Ɖ� eX��v��B-�?>��IQ}��Х�,m_����銾4��GĎOa*{�lH�*�{P�WVȠ!�V�C֓�n�A�pf��G�J��Q�p����1"i���Hm7�B�岅�J��p�d2�=��ܱ�7B�x(a{f!�KH��ݠ.��e� C5̒����!�b�f�� �{�w/��V��8����b�A�ms�����(,��S��?�UK�P>�?V�?�w��0����D���Fo���
��^�A�AM�կ5�Pw>�|Vj�}�jx�����w�8`�ճ��iޟ�v_��zC���AĴ(UW�/ە���S��uQpdX<�L8���͐�2(��	^}�V�E��-�@:�h�ib�@�>����?9�'�WN�	�'�*2yE�Y2�R������߆���M�x^��4���Jy���z������)�@�� Z�>�I;v0Q���UaF��G�h5����;^��Iy(����tA����,�p�v���d|�����Sz��`�6,��Z\�A��W�Z�"U\���9_đO�6�H��|L�rK�%׆$+'�� �C�l:�d��M>[MP��t$Á���b����N��|=13~������R�e�[��0�Q�E�+�����i��c�Y�(s�|���;)���6.U����Q\)�7���]�������r�K�U-�a����d�M5Ϭe�c2/~'�Mt�t���M�E|f�)�c���ů�g��-[��TK���o&frN�(�m���8��\g�ֵ��NE�=P�R��v� �sP�0ЅvF�8k�-��6�k)������\��3���K�Uϗ����܆�Q�q����f�fܿ��j_!s-}�_��l���tBNzC�n�>m'N
>�?@lLښ/���.G�z�d�[]1��櫍���WJ��i�(�=b.���ԭ�cjܡ����&�d�'�����>��+Y� #���j ,ʹ��k/E-���`N}Lk'��bn����z~[��'�c�qD�����9Ӽ�Q$���}f������*x�ГA�߰��`߂B�AY�9c���Mկ�!���j�n�9��Ջ�F> �x���!��X{�am\�'�cuה1P��-�=:�˭Q�z�����fp��τ1���;�f��C!C��?�����Qp�®6v����#�|�d`���*�ׄ�IW�%*�Q��"��C�CS���ÊXí DNT76w�B��O3���- �J;w"o�M��p�}�C�Cγ���h9
JQ�Q����QQ�(�zK{�н���s|��J��