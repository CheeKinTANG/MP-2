XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��KP����T�����Os�#_�ĀU�Pw)j�#RT��n ۈ'��{��s���5�G�%�3��@����^���
F���&I�<�Gh������fhdU��RR q���m�Z�po�H�9F�3���Y�=��w���c���:~�Q���E	�eu�uW�ܹ"�C�sUb5S�n&d5K'7�������ԁ;b��/^�j�����}�覩���P�[uf�-��F�I�н-8�����U8���)g�8�M�k��3��M�ew�R��`�D�-��A��(��T1U���w�����\b7�M�B�4�}9�	P�%
+p ��^�����O�[��Q�UQ�^X6㔸�7�@���u�s�H�$M��@�wvc�i�����s�����O"9KSZ{E��Qr3~/9NQ���92a��V��Y�.�Ywր�!����T.��/v���2R�����Fk�Xp�@���L�p�Qx���ń� ��c�Yv����j<׸���ޓ�]�!�&� �y�۶��z�S��Tu}�I|��瘨��+�L���5�m���YlR��4m$��>�XPf�-K�wRX����[<5��@OJ��nΈ�W��0�Ғ�6����Pؓ���"8�3�J{���Nw��q�o2]s����a[�K4I%g��p'�6[X��+����ޯ����*��c���󽨇���dM��V��"z�m�T畘p����9{�%���
�q��z���*t�a�Q�������j���XlxVHYEB    3b09     f80#�<�u��,�y��ܑt��ԛ��q��r�H^�U,"&*�e]�P�g�RKF���q&�"��p��V����i�c��Y�,4Pf�i�����	��Fj����'"�����J��4z�8�q�^�?){r���9	G��� O����<��&�l�;�<�h6g6@X��Z�@��8Qy��<^�7-$��l��]�_�VKx���9ܯ����[��W#�6�O�~�&����Zk�}b]]�=�0��!�8|�I��h�����Ηa�/�����MwHGhlq����o������7��m\�Z��܌�G��R(.� 'R.� ��0o��P��}B�a����8ZX�"�sS��9��������&��93���řҳ`߄d��� A8�]��|�7E�<0^*��� מjg�>}���FS�lR����t��,���@���aЩ���q���@�GF���2�=���!Ja��k��58ˤ�9�٠�|�19ynE-��ΕO(�N�a[�z�!_�r�$�����1?�%h�c����f�R���0m�`Y��סFRME�Ǳ�����.�8���xBSX&��,0N+� ��զDB��T��E�`��k�k���'���N|q1f�����v��w>��m�'!�#L4���xfG�h��tse�#ڙ�D�R�Y?���.?㎚)\zoD3Du�5��UTC�w�J�J���oDV>�"n��;r$|;?J{�����N�c�=h��:I���QV�zqgY���K4w�G�� 8�{�?3䕜ެ���[�BC��^4"�_k��aE��D�M��F<S���V��ĺ�^����KM�y�#u)k7ސ%Ҫ=/w�(����3��ƻ���d.9�k^ɷ�	N�\7ࣵ���?4��'2]�R����~;��@A�!o��S�A���O x ��(��y��gP��c���֭_į�&��Z^��Ȟ�����/%��Y����SJ�;bR���� ��V�0�����Z_�+�e�\6F��#E����ܮw`|��}k�.ױp\ҍ^�S���v�9,�oW�d����X��r�uHc:{$��?�� +Mkk|��NF���
��l��E��'+��Ҫ2E 1tb�0?��g\�w73|�]���^`���M���k0h�kI|z��T9�^K2����/|;ߥ�0!zȘ��D���Ì�;������e���7[�0�ϓ���}�H+]`M�R�7fd��D�r\�Q�}>P_�p7ިȗ����㻧��cS��h�,����Oh�'��۹���Œw3�F!l�&��3M����.Ů �(����v��%ak�ui�ڶ[�9"��+\�@䏃4�!�T�-��g�U�%�ޙ&�e���i��|R}S]s�
*f� �F����پYh�Z�W͛��{�D�
��'��\�HP~�_;;����NI���_K���p�:�����'��D�9ߋ����G��f���A5�{o�L.���?�m~���͍��4��(.[��V�����tO�#j������'������w/�z�V�_.��@��������]9��1�9d[���z���t����)睻{�h�.3K$&��W;d���R����'�'��I�~ݦ$l�{V�e̛�k�T�~!��U�xϒ�(��f��xr�H�J�I�6��|w��?����VieS�y#7�޼y�CG�W<��tO��s��� -�������k�Q[>5{x�H�I$�D�Ӆ�35�$f����r�cLV�D�#0BJ۶!  $ɿ�>�VS- ��3�D��KºY]cq+Q����Q&�!? ��9��������sj��5��i{Q��}�����0hPQ���^J���P�3|כּ��K-�����6�)�-��X�|��H�-���[�>�?j�{��Գ:�͚�:��j����a#�c󕢦m�	I��}�WqY:���'�|�?#*Z��g,X�$H0����Klw�C�O���uK^j�}6�/�.��EY��!��f���4,m��{�:l}0��vy��Y+��a��� ī�Cm?�Z�;(��SU���t�"�8�~�ȧ��?��R5F6_8-a��[�z�@C�|g4�&�uey|j���y�!\��I��D�)@S�cj�n��,����kw�d�q��/!/�ԁ$zR�&L�e�bd�.�p�Wz@����̨��}�U�(�;���Qaxo�PԿ����NV�[�֨ƥ�j,��k�9o�����m�eҶT���Z�<��/J�p��!�5�ɞ�¨��?��y���}^�P ���9~�Y��t%�U)mx����%o�������:*��������o�:�hK�<������6�9�~	�=��JsqxKF�ШJ��S���j��7���ʧ?ӿ�蘲K=����~�]�S��<¢g�B�%����$����G?RG֦��p�SDo+$���Ui#�Ϳè��\�0Tn�ט4��0t�&��T�ݙ�'v�m�{N�+pä�Z���$4ߥ��n�a�ًAiA���0���)wiƽ�)�,����T�eS����Q{^(���G�+0�sM�<�ɐ�����tK��ꎪ6?کo�&Tv��-H�H����)|az<o��l�c�R��/�-�]�T�̲%u1z�#�䏟�v5��^��MfM�N�)��v���o�y�E�Q�v�U,E:R~꒻�W!����֕��!aµ�,i>I�1�O�׷�ThX%]`a�����%���M����P��+�R�	 �[8J4�Ѓ�-��1�7�. ԃ��Tc������c<D���P�b����)�����f��Q �Ү:�?7�I1������Ӄi�&�K	ϐ-V�M�-��Z���~5��6}LV\����:��57�}���Τ�(�+V�+ ���d:�e�����W%���q��h5;��>�Q*F���92bb�����/��G96$�K���p"������,�2�3�C�P��}�'����Q��]����2���³zUI��I�f"Mӆ��]�؋*�σ��&�fj.s��¸�O6��QCT�.Ϥ�Z�_��1,,p߲�T�̃�n����:��p,CC�ʞ�k0Ty��=��Q\.c�kZƼo��k����t����4B� �=o�Y	���]}�Y1���#map�psR��pQ�,ng�;(�H��"����b9��8@�RJfIhA�Wv��+)qJ���AF�j��]o���Н3Gd�D(�n�ìΣ?�^uC� Jw��O�
��R��.H��fEn-�����/d���Sc�vg�Ċ������JϘ$�W[�&'8ɡP�t^�s�i}���U�\"��5��0�e!���\@�N<j����%�����p����z�`�J�bm���W���kl��,
��B����xZus�E���c΀���|�������}�_a=0��Y�;K�װ���}q��fĚ�2���L&B]���	`5϶]d���[C��/��߹����M��c�}8F�]��lW�aF�/��nݩ�8��q�ؠ>v�o=�xG��e�51�/���säK�99!;if�r��},|�cs�o�������\�fF�H�^vJ��<���ԇNg
.s�ѯ�3aM��^E��NtfM3���0�I�������AXFJ���̋e�i�ݙ��.G��K����^���$聹M�w�PN�AT���ځ���HJ��`*6��#�*�P%J~�ɷw�D�>����B��^���u��o�cl0A9n���!�'b��B��Ƨ�t71"���	��7]�v�<�K�3QDasL�O����/��#�BÒ�u_h١��I�@z��u͆��N}�����8