XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��½oB�KI~���A�1F����r���Y7��T飫�w��H�  f'׼*�o��9�)�"5���";]�_1�Ex��+8�޹�|}V�����豾Yiw������Ǘs��;P{f&�As����X\��z1�"ŌH�J�V��/�=��#�z�TG�oR�&�����<�:y�
�C�X��Ř*��Ŭ+_�ʢ&
@E�G4�����9^-rp�m�۲;��ɟnm�+��8�X��uc� a�.�����3�۟�\��mgӽ� �D�WN�g�Jص��M�H�F|\3���:j���)��v���ӓ��;"*�Ŏ�V㺨[Bt��['�˛�xg�遞�d�\�*�T�A\�8l�q>Y���SY��������kF�
m�L��R�Ҵ&%l�r�(=���7��-ЍFd��N�[�49�-\~-�Q5E�̱h^|)#�������x��mV�b<{ኼn����'M7�s�1��'�^�3(q��_�BoHm-5&$,��������?�-��G3r��#��:BK��4uQ��T�n�I��
�+J�64V��#B��{-���s^ �4I�s��1������Mq���G�ͺ�9��>BN�-f���탽8ep���*�Y���{�>A��h����v�oJ�5lx�y��Gfd����������,�K���Å��G&�.1��:�����[	;��{_���0:�"`t�N���ykЯ��.Y V=��g����m���XlxVHYEB    4284    1110�����G��#�o6�Bمj���SV���w���B���T��'���?V��b���Z������,�J��@��k��.��{�~(��8avj��
)�<"��/��I������n�[������0t���<Z:F^�q=3u=�I��V���B�Z.�����
l�zfJ��\z�Z͒�&90ZI�<�dL���>�}�D���w�(��;���%��3&з����6�-\9BX��y��\�ޔ3��<��"<^�J^�b�^ r�ҷ߬��t�2l�κ?���_�?m1�o�beS�����|���D(G�-7�9��B�@�u�0�	W�+lppXñ�� �m�� �q�<��;�ĭ�/����x��fH<FՎ�n����7��W�1�t�sr�����: :�auGHl7e̍�|�XK��0�v��f��[��7���Cۄ�$SZd�O��8p\�w�j=x�tU�Q��1�&�M�@�χ�6ҳ�����/6�ߠ���߳�z}�Ic�D���v�I!@����k���e�>%�Р(��6a�Bd��Ap'aֈ�XH��e)y�_�^�,��Q`�H���5FyU>[�!��W<P�2+�82�H��~��q�D3|�$���C���[��'U���9�?��ڗ���Ÿ��Z|�u���\�\�����u2
1٪��DV�[�j��)ٮC_�P�F�a|���5X�W�x��H��Fut�wb 	dR����xX"KK�i@W�����͇�������^TD�pQ7�׬?$�m���{!>x@Jv#��uv��y�k\ EYV٢7�+�(Ą��h&��;vP�G9�iJ���^�j��G�M}��c6_���(�����A��D2-�p�=��rǥ�@SE�#� ���Ê�~����8�N{�J\T��s�H�5zD�Z���ܕ ��z?����K�A�i�3j�&ΐ��g���Wf��G��R�c���d�vaMO\6^)c�J8���_ML��o��-%s8�U���R�q@�����@K$�X6�v��5��<���	J_S<��?�t1$R�V��N�����������v"H�g�}�D�ݲ���*��Ć��{6 ���X�8���e,$pT�L^T�R]|*���v��o=�`uJҒ��X���0�� ]f����2b�[0��}n׿zM�l��(G���h�1�+���ZX���[�R/�Xo8:��(��|��sc�aZ�%��l��K��i��1�����ofl/�l�b�)�!�癨P��B%���p�`�P?WTt� i}�B�yV�R���a�`����焱�z��}5M�O9���r<�l�����ؖ�6��M=aG|N�@�qj��_���-g�&v������-i�n��M���'d6�ɋ\���H�V�R�N�-�G������|���\��֥Ȓ�s�&_����|rrhJ[��d�靯�MY*!��kH�Vz�6d�)�<&ݟ���x<I�W�k���ղ�0;U�.k���xe<�l��C?x�#B��W��r�P��e�vr�c�e��4�6���3"����3��ۀh�@����xi���+	��F"�.����Ė`����ul�p�n�8s�4Q��D���[s�o���@lc�QJ��]I;�m?&m}2�	�7��.�8�#8��:s|��u��!F(P��ޥt��$H�V�
Pm 	�'ap��I��)��h��"@K<�1�d�C� �װX^�%��Ϛ]^aj�靲t�h1��e���:W_���ʘu�]0��*Qn�˙�$����Y)�����DFҸ`�'&<�z�eh���~��ͨ���#7�L�걞�?P1�����S?#X��4q��T8U��7����Ob̃o��(	`ͺ�1�P`f��P�Ƶ���ч�1��G������:�Rb��Z"�	�:�š���Pؽ��x��������'��	���l���0$�3{�!�l`������&]�L����{Vg�����_�v���S��̕\����h�D�kߥc����;��9�W2��u��x�|5��%M�{I"h�}C
@`+N�iD���� �	�_�5�^`G���/�9���H�;��uӒ�����N�.��U0b�/$�DL�SF����<h�OpT�pJd@�����p��`;���yGUN v	�ռ��m��ʇ�K�i��(���7g�_���gE6_�!�H�|W/^E��*J���R�<Q�!q��.�rK,�!̣V��J�w4���E�N�9�0[i;*�����2gwz�R>���c��e �����ɱ����n��X����� /(�Z�1􌤍[��3 F��V0��
��)��i�+1;��=:�h�����lLIe�|x��5�f?��ۤ���H�N;`xw�
TZϟ�әP�B ^w`��ۀ%8�/%n���y�jt-Wf �\p���%ƭ��y;�Ln��g��A��Y��c�҆rn�`��P�cdy& I��-�m���M��]X��0���Y�K&'Zԭ {ګ�4|Hi�wG��Q�J����QA@��攁>�YM����^�a�b�u�.g���uRk�}jv��<���z����c�Ja�t(ǾF#Ds �X��_���n�4.���i1�}≧��N1s�<Hގ"�'-L�#��+��u)�����b��,�q='�x�?�L�,�{&ٍ��q��n^Q�"'qPC��D�	Q���������q@��.5�%_�=�ڴn)�BX_ͮ����b��C'r���/��ZX�5�S��xy���`�)�����Y���'��g�N���%�������}�����!��OS%i��넮IBY�w��>,�Ա����Y�/ڌ�t�؄w�0I���`�r���4��Fդ"n8�����A1�4K\X&�&ny�H��E!��`�=������5�V���-ό���S����+�ť0q*R�� wFL�y�2=�1��97�l���/1�|$�-�4 cgy�!� �aq'�v�Ѫ�ԍuÁ�Ғ�Q���K�[�:���6�8&�ޓ
�si��[|�a�Z ����P��s��I�c�@����wԀ¶���J�y9���y���@�ĴUm/ße�?�*��9��@��CTR�����}YMaF~��O�g!{�V3$�X�]�C�g'S\J�I�(=Ҷ�F����4H���5W�n�_�|�c��9��;��9�g6D��P�����MJ2��`��DF��$t�,���l��k�pV�����_�5Gc~pV�kVހ�
�^���,��B�����-��$�����	M��m,j?�ܜZ
�s��62��`�y���'�h�G��aс�rKG7j^s�J����@�R8Zh��(� ;��߀��iJS��r���R����g�Z%ٚ��G��C����?���x��X:Ko*�,�E�����p�Si˷Ӣ�A/��d����;t\@}���Fϛũ^�ٹ|t�T�28N{���R����^�$�=06�̋p#���z�Ѓ�R�k��3���dSQ���7��?=O�^����ւ^F�/T�$�vm�,;%+�խ�B��!Wk��鐌�����1>Yj�����b��5�n���P3K����&�N�0<�Ze�zʗ	I&�r����,n�F0��Z�]n�XVK���8е3��i���7���PU�%E-juV~Vb#c�c������TYY��lh�z��?3S9ł��.�#1��(�S��?���"��C�&qo�$��I	�b�x�����f��i�l��?ȚٯR5�����ٹ��a�} qA������ �,�趥�����[<��b�!�Y����"kvЮc>�W,B΃B�{��e�3E=A��N����n��<-y����O(tmI����W<Q�tv��I�y����\L����)Y��|U�gf�Ʀe�����'�S�:��.Uc����d�4T�L�`�.���n8N�,x7Q�6L!�}O?���p����y ���"�5򜣮�G<�$��<,L��s�j(�HS�}�h�]sM��,(�TT�k��E4A����e�ŗ�(���7��s(K���ӟ谯���֯~�ǧە�?�-�Ӓ1�$N�f�F��'�Y�.���b(ٮw]���Ȍ�0�aM�4�Db;T�S"����{X?�:��˂*���dd:	"$�Ք�
�Ūj�e6W����^M�@1�N���(&di�g�,�iU�	*'^5^i���B�Z�����T�$��Qc�A�X:��s<