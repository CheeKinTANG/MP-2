XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\̛&���w(���R�a
����س~^�[_�|�b;t�b�Nf
�J�=�|��^ҋ+�.��ߓ���eZz#����+4�k+_���:x��B	S*F��^z�;HwD�\_�g��QQp��աK�	J�p����"*�#p�4
�8�v���j�]ޖ�#@���~ ,?�D�l1�P�&����?yqք��pK��z�c���1���i�g�+���S�A+w��)W�Q0#�ϴ+j@t��l�` ͽ���Y[ �Z>_z�2���|ݼ��C��8��O���U5�LT�q�O�5$�!C�Bl�8�g���^E��j ������c��R; ���^�ωwC����TȚ	��;V���T]v� n�NLg�'��� ���Y_a��[_$�Tw��"�p֜��e�@dt��r�tr�ǵ���arc�l4n��4�6����[�cn���N�������Z@��/^�O�MC��YE����uބ���pk�^�5����7:���C��|Q��W�y��X|(�D��?�ҵ�dn2#t���"�S)i���@�k���j��wIw�G6�HL6�~M�]]��%�)� u���E:7�Q��F����Bљr*1�fv�T��\��Q�fs-��B�=4C�ͽX�frg������1t��JD�w4`n�#��Et��]��~!{+��K1x����ۖø��L�ms8����v5$�� ��L���ao��绪x���Y���{I��0[���N�LÞ�g�$XlxVHYEB    4284    11107A�v������Ǐ�a���Xܶ�Y��Yd.�w�=��ީ��X�<��/R��gF6�}"�Q]��m�E�6�U2�E�Y粹��xX�jă|�Չ�pCN�3� n��7c Φ[Z�VÄE�=����e� j�.A�1^��l�*ӈh<1�Q*.�s:��c����Q�?C�z�,�(��<��h�[��*���#V����4C�� !sD�D�1�7o}"��틦v!i��P�5V*|���߹���d�󷳶F�t� _��e�T@+������� K�4�&�_c��"�II���57�~o�R�a�T�D7�C���S�<qo�x���0㳕L�F����"���s���w)��pߨ��|1�s̀��@��ǤqeZ���}���q:μr8�s��Z���u���jѡ���(�6BB±nVk��Hez�$3gs쭱auw^�&<,%x=�&��n�#�u���%�+J��ߙg@�g�o�9cx�c$4����?j=~QsU�H΢�����ɼߗ	�~Yr>#���� ߔ�vZƫ�5D�R��Ҙ���f�І+���E�X/H�R؝ũAX��<�i���z:�x5X�a����K{9�>#�� �,�����G�y=����EZ �n��|]�Q+5u����7�x�\*@BI���f���n�ї��t���p�G�6��ܢ��o?������3w&<`c&E�G����/�O�J\�N��4��	z�k��o�_����}!r��f��W�$�:p�z�M�M���\ �DqGQ-�W��xVw����'ph�P5�R ���>���RP��,�J�L�Q�^zj���FëH��VBSK��{�U�����0f��.�[
&�[L�&N"�.Ǟ'}4��BKX���A~��Z����O��÷���B/8b�1�mg�k�p�x'�����i���.	�
�`P�E$�n��r���;K�u!�N�8�<�:�T3����B�L�@�/Tg*�����h�� ��	��޽����D�#>�A	"sȻ>9M�	T���@�q#k�7Y/�nOV&.��4�˫ww]��u�}њ']�}h0����Χ����K}a��Y���S����>�"!������~��{@�#��R�&���k�����W(�[�-�c�h~3d}���%0�/�\�ӅH6�]^{��P׸�{�u�M<�ݻ��}���>s��ۂ�Z��eE�doUF፵D��DN�}<��dq<Ftd�����M��*`����=��ךI�&��'���w���Hd��߁pCO5ע��Ґ��S����s�%s�T|v���:�2ps��-���6ju~�zn���K�1� �F�c����?q��T�7�^��:ɛi�>�W5fU�b:X���̝̅Z�m��$?�#��A���4S�Z��驩B5^��1�V��Y��G�I'��M�xq5�)y��Dk	��ŉw�.�]ETueQS
5��_i�/�,�qU��+ؠ,�Ŀ�<�(��P/�M��-�v㔠��Py:m��h����q$�U�X�;U�� ���1��Z�7�ZUE�hތO�qMP4F���S���!�]�b]�	�ym;�AF䣦{�om=�����o����/Xh�5L;n0���a}z+��*�O��O�]u��._����)��ZK>���q&��}�ݎ�s�K���j��R�k�%1���A�<�Jӹ Q�j\�P'��/|Ф�: ��I�rJ�n�C��y��k�)�F�SÜ�fY���c�v��q(ՖBk��H���l�sR*�.�e���G�Wѱ�4:�@�婆p_wboR�M����
�M�����R�
�sw~]q���4w)�����Q�Dwr�.��W|1����`GtX��K#��~��Z{��n�_��gI���'{����@oٿLY2v`���'�}���;��-���A�����}�`_y�U\��<�@-��\�������{�8�7�H�<rPz�%Ka�g�c� Z�!�əl�W�V� $(��!?�"��>S�$I廵Y� ?�Bڧ~*��~%�0�~��\�~նm��%��|c4�S_'��&k�կT[��p;�G�zG4RxVw��gn��L����ռչ��Mŷ�n���W���$�$��4���u�݌B|̈�\˂Z�J��<(�Y��G�祗�wp����]2F�����44�V�l9@�e��&�[^�/Fy�:+�^ቋ�<|��jF7@��CE��2��X��C�2Yb���S���1�T�
�ƣPE�c�2�n/�q�ı��;<����Nra��xR��)SHp�@�3>�@=�v0��oȲ=���/ɤU�TRx� ��E{AiB����7����zy����eMGU�Z��u$M��AR�1��˛�����ْ:�z��b��~H�.9�B�_�:hH!,���a��
=$���vʉ�3[��GZ��Q�@��=|,�-��V�T�&:���W�=J�l�hq�Bz��I��2�A�D ^$�7�ܺ�+�^q�/]3�Y�z���ui�us���ƅ��gL%�ܮ:m�G��Д���E����v���;~����h �9�ڲ]�'�;=H�U_`U���v4{�0�?���@�R�vz� ��\��74��@��`���ٯ!�Q�f�r���k��`y���=�2Vr4���m��Y[ )�d�/FE�bB�f��'��C¡\*����{��Y�Y�u���>5��X�v6+ ה!b����JZ�hl�~�hvc���baI�q'x�D�.�֫ ⎻����"�����UHwh�����/���-(a�����ɓš�*��r{C&H������[��=6��������!�I���5&n����B�u��O�n�=E�cE[��Oz/�5jq��h�*����m/��H���b<�W����~��7������!+�L��M�����ǁ*ꖣ>��Hɓb3�[o���#%����3j�\��J'�1���΋����kG@O���g�j����dYH��M�W��u(MT��
�*'�~���E�=�$���n�p�8{?!\�'�v?�i�&�
o����\��z�6��y�.sE�/}�:��Y�7~�<v�1� ���RB�U�+V,�P��L�hk�>Q������YN�HX����g�>�z���an��$���V�LO�i��JMT]!)n�t�� #Hd�x�\����2[��E@�/_Y%۝�׶��<9�������v|������[�R, K]|(
8�Eˆ�I!`�}��+�@�>C�+�,�釂�fOg��w�~u.�dE��}?�iqQ��Z������Hiׂnx�w��>k�-7�%����2Yj�-�׽���#$����cA��Ƴ�Ќi�f�?�"=[���m? r~_q�J�D���P���ق޺)��_�*]F~���3��j��qo:�*-�d�Gh�a:v/���B����>)t�!pH��J���U?bEs����?��E˒ADֈ����1�_a��i�@?�c*���xIp�\��Y����d�:R���H�	���K]c�J��{���B�!2ȣ�ch���F���~�JHjX�t�S�4�8��3�%�T�j����[�*9ؚ5�y*��}��������#�y��33c���{������'͏os���M�P'�ȩt�^���1��U�~Q���k�|��o�fg9_��ϴz?��ͽoq7�1����l��qF�o%��]�s��I�qn��q����"�*Rl�I�1�L�U��cf����E#�*�EO���IN������o٦��h,��e방�~�c�޻��hH� ������l/	�WX�,�C�L���� ���,~Xr#�����V�7�]�7��b(4QH��d���#�1��:-�X�/rU��D��f�k@g��{J��Ae���!�-p��X�g����I|?-�i<+��*Z�rZ���ph)sm��Sk��6�H��J�lB
F0z����L��i)%ʐܴH��u��d�����p�v�9�ٝ��Om6�3��� �
GG"6�k��%G�	T}�7��ID��z_Q3���"��f�X �Rv;�7�I�!8.	��=ր��fX~W$��zs�/�_z-P��YL֞���Ю�+�,+]��L��kc́9��7��m	5t?�Բm�|��k�t=,E������.����&B?5Y�1y�/tJ�.L�~�U��X��Hq'�8]��,�kr���A